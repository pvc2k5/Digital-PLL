VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

VIA ring_osc2x13_via1_2_8960_1800_1_4_1240_1240
  VIARULE Via1_GEN_HH ;
  CUTSIZE 0.26 0.26 ;
  LAYERS Metal1 Via1 Metal2 ;
  CUTSPACING 0.36 0.36 ;
  ENCLOSURE 0.06 0.32 0.01 0.06 ;
  ROWCOL 1 4 ;
END ring_osc2x13_via1_2_8960_1800_1_4_1240_1240

VIA ring_osc2x13_via2_3_8960_560_1_8_1040_1040
  VIARULE Via2_GEN_HH ;
  CUTSIZE 0.26 0.26 ;
  LAYERS Metal2 Via2 Metal3 ;
  CUTSPACING 0.26 0.26 ;
  ENCLOSURE 0.01 0.06 0.06 0.01 ;
  ROWCOL 1 8 ;
END ring_osc2x13_via2_3_8960_560_1_8_1040_1040

VIA ring_osc2x13_via3_4_8960_560_1_8_1040_1040
  VIARULE Via3_GEN_HH ;
  CUTSIZE 0.26 0.26 ;
  LAYERS Metal3 Via3 Metal4 ;
  CUTSPACING 0.26 0.26 ;
  ENCLOSURE 0.06 0.01 0.29 0.06 ;
  ROWCOL 1 8 ;
END ring_osc2x13_via3_4_8960_560_1_8_1040_1040

MACRO ring_osc2x13
  FOREIGN ring_osc2x13 0 0 ;
  CLASS BLOCK ;
  SIZE 126.285 BY 126.285 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER Metal4 ;
        RECT  117.04 7.39 121.52 118.05 ;
        RECT  72.24 7.39 76.72 118.05 ;
        RECT  27.44 7.39 31.92 118.05 ;
      LAYER Metal1 ;
        RECT  2.24 117.15 123.76 118.05 ;
        RECT  2.24 109.31 123.76 110.21 ;
        RECT  2.24 101.47 123.76 102.37 ;
        RECT  2.24 93.63 123.76 94.53 ;
        RECT  2.24 85.79 123.76 86.69 ;
        RECT  2.24 77.95 123.76 78.85 ;
        RECT  2.24 70.11 123.76 71.01 ;
        RECT  2.24 62.27 123.76 63.17 ;
        RECT  2.24 54.43 123.76 55.33 ;
        RECT  2.24 46.59 123.76 47.49 ;
        RECT  2.24 38.75 123.76 39.65 ;
        RECT  2.24 30.91 123.76 31.81 ;
        RECT  2.24 23.07 123.76 23.97 ;
        RECT  2.24 15.23 123.76 16.13 ;
        RECT  2.24 7.39 123.76 8.29 ;
      VIA 119.28 117.6 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 117.6 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 117.6 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 109.76 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 109.76 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 109.76 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 101.92 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 101.92 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 101.92 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 94.08 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 94.08 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 94.08 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 86.24 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 86.24 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 86.24 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 78.4 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 78.4 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 78.4 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 70.56 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 70.56 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 70.56 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 62.72 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 62.72 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 62.72 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 54.88 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 54.88 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 54.88 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 47.04 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 47.04 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 47.04 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 39.2 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 39.2 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 39.2 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 31.36 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 31.36 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 31.36 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 23.52 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 23.52 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 23.52 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 15.68 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 15.68 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 15.68 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 7.84 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 7.84 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 7.84 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 117.6 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 117.6 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 117.6 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 109.76 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 109.76 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 109.76 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 101.92 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 101.92 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 101.92 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 94.08 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 94.08 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 94.08 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 86.24 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 86.24 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 86.24 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 78.4 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 78.4 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 78.4 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 70.56 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 70.56 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 70.56 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 62.72 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 62.72 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 62.72 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 54.88 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 54.88 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 54.88 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 47.04 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 47.04 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 47.04 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 39.2 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 39.2 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 39.2 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 31.36 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 31.36 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 31.36 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 23.52 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 23.52 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 23.52 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 15.68 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 15.68 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 15.68 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 7.84 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 7.84 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 7.84 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 117.6 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 117.6 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 117.6 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 109.76 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 109.76 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 109.76 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 101.92 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 101.92 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 101.92 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 94.08 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 94.08 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 94.08 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 86.24 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 86.24 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 86.24 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 78.4 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 78.4 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 78.4 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 70.56 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 70.56 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 70.56 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 62.72 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 62.72 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 62.72 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 54.88 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 54.88 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 54.88 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 47.04 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 47.04 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 47.04 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 39.2 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 39.2 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 39.2 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 31.36 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 31.36 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 31.36 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 23.52 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 23.52 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 23.52 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 15.68 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 15.68 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 15.68 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 7.84 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 7.84 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 7.84 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER Metal4 ;
        RECT  112 3.47 116.48 121.97 ;
        RECT  67.2 3.47 71.68 121.97 ;
        RECT  22.4 3.47 26.88 121.97 ;
      LAYER Metal1 ;
        RECT  2.24 121.07 123.76 121.97 ;
        RECT  2.24 113.23 123.76 114.13 ;
        RECT  2.24 105.39 123.76 106.29 ;
        RECT  2.24 97.55 123.76 98.45 ;
        RECT  2.24 89.71 123.76 90.61 ;
        RECT  2.24 81.87 123.76 82.77 ;
        RECT  2.24 74.03 123.76 74.93 ;
        RECT  2.24 66.19 123.76 67.09 ;
        RECT  2.24 58.35 123.76 59.25 ;
        RECT  2.24 50.51 123.76 51.41 ;
        RECT  2.24 42.67 123.76 43.57 ;
        RECT  2.24 34.83 123.76 35.73 ;
        RECT  2.24 26.99 123.76 27.89 ;
        RECT  2.24 19.15 123.76 20.05 ;
        RECT  2.24 11.31 123.76 12.21 ;
        RECT  2.24 3.47 123.76 4.37 ;
      VIA 114.24 121.52 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 121.52 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 121.52 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 113.68 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 113.68 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 113.68 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 105.84 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 105.84 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 105.84 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 98 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 98 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 98 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 90.16 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 90.16 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 90.16 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 82.32 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 82.32 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 82.32 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 74.48 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 74.48 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 74.48 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 66.64 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 66.64 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 66.64 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 58.8 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 58.8 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 58.8 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 50.96 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 50.96 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 50.96 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 43.12 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 43.12 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 43.12 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 35.28 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 35.28 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 35.28 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 27.44 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 27.44 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 27.44 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 19.6 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 19.6 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 19.6 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 11.76 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 11.76 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 11.76 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 3.92 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 3.92 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 3.92 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 121.52 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 121.52 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 121.52 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 113.68 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 113.68 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 113.68 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 105.84 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 105.84 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 105.84 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 98 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 98 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 98 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 90.16 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 90.16 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 90.16 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 82.32 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 82.32 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 82.32 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 74.48 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 74.48 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 74.48 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 66.64 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 66.64 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 66.64 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 58.8 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 58.8 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 58.8 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 50.96 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 50.96 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 50.96 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 43.12 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 43.12 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 43.12 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 35.28 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 35.28 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 35.28 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 27.44 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 27.44 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 27.44 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 19.6 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 19.6 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 19.6 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 11.76 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 11.76 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 11.76 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 3.92 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 3.92 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 3.92 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 121.52 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 121.52 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 121.52 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 113.68 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 113.68 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 113.68 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 105.84 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 105.84 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 105.84 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 98 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 98 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 98 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 90.16 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 90.16 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 90.16 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 82.32 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 82.32 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 82.32 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 74.48 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 74.48 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 74.48 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 66.64 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 66.64 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 66.64 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 58.8 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 58.8 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 58.8 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 50.96 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 50.96 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 50.96 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 43.12 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 43.12 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 43.12 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 35.28 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 35.28 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 35.28 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 27.44 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 27.44 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 27.44 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 19.6 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 19.6 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 19.6 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 11.76 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 11.76 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 11.76 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 3.92 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 3.92 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 3.92 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
    END
  END VSS
  PIN clockp[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  87.78 125.765 88.06 126.285 ;
    END
  END clockp[0]
  PIN clockp[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  72.1 125.765 72.38 126.285 ;
    END
  END clockp[1]
  PIN dco
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  124.74 125.765 125.02 126.285 ;
    END
  END dco
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  77.7 125.765 77.98 126.285 ;
    END
  END enable
  PIN ext_trim_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  123.62 125.765 123.9 126.285 ;
    END
  END ext_trim_0
  PIN ext_trim_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  122.5 125.765 122.78 126.285 ;
    END
  END ext_trim_1
  PIN ext_trim_10
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  121.38 125.765 121.66 126.285 ;
    END
  END ext_trim_10
  PIN ext_trim_11
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  120.26 125.765 120.54 126.285 ;
    END
  END ext_trim_11
  PIN ext_trim_12
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  119.14 125.765 119.42 126.285 ;
    END
  END ext_trim_12
  PIN ext_trim_13
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  118.02 125.765 118.3 126.285 ;
    END
  END ext_trim_13
  PIN ext_trim_14
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  116.9 125.765 117.18 126.285 ;
    END
  END ext_trim_14
  PIN ext_trim_15
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  115.78 125.765 116.06 126.285 ;
    END
  END ext_trim_15
  PIN ext_trim_16
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  114.66 125.765 114.94 126.285 ;
    END
  END ext_trim_16
  PIN ext_trim_17
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  113.54 125.765 113.82 126.285 ;
    END
  END ext_trim_17
  PIN ext_trim_18
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  112.42 125.765 112.7 126.285 ;
    END
  END ext_trim_18
  PIN ext_trim_19
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  111.3 125.765 111.58 126.285 ;
    END
  END ext_trim_19
  PIN ext_trim_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  110.18 125.765 110.46 126.285 ;
    END
  END ext_trim_2
  PIN ext_trim_20
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  109.06 125.765 109.34 126.285 ;
    END
  END ext_trim_20
  PIN ext_trim_21
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  107.94 125.765 108.22 126.285 ;
    END
  END ext_trim_21
  PIN ext_trim_22
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  106.82 125.765 107.1 126.285 ;
    END
  END ext_trim_22
  PIN ext_trim_23
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  105.7 125.765 105.98 126.285 ;
    END
  END ext_trim_23
  PIN ext_trim_24
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  104.58 125.765 104.86 126.285 ;
    END
  END ext_trim_24
  PIN ext_trim_25
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  103.46 125.765 103.74 126.285 ;
    END
  END ext_trim_25
  PIN ext_trim_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  102.34 125.765 102.62 126.285 ;
    END
  END ext_trim_3
  PIN ext_trim_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  101.22 125.765 101.5 126.285 ;
    END
  END ext_trim_4
  PIN ext_trim_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  100.1 125.765 100.38 126.285 ;
    END
  END ext_trim_5
  PIN ext_trim_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  98.98 125.765 99.26 126.285 ;
    END
  END ext_trim_6
  PIN ext_trim_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  97.86 125.765 98.14 126.285 ;
    END
  END ext_trim_7
  PIN ext_trim_8
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  96.74 125.765 97.02 126.285 ;
    END
  END ext_trim_8
  PIN ext_trim_9
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  95.62 125.765 95.9 126.285 ;
    END
  END ext_trim_9
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  78.82 125.765 79.1 126.285 ;
    END
  END reset
  PIN trim_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  94.5 125.765 94.78 126.285 ;
    END
  END trim_0
  PIN trim_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  93.38 125.765 93.66 126.285 ;
    END
  END trim_1
  PIN trim_10
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  92.26 125.765 92.54 126.285 ;
    END
  END trim_10
  PIN trim_11
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  91.14 125.765 91.42 126.285 ;
    END
  END trim_11
  PIN trim_12
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  90.02 125.765 90.3 126.285 ;
    END
  END trim_12
  PIN trim_13
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  88.9 125.765 89.18 126.285 ;
    END
  END trim_13
  PIN trim_14
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  86.66 125.765 86.94 126.285 ;
    END
  END trim_14
  PIN trim_15
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  85.54 125.765 85.82 126.285 ;
    END
  END trim_15
  PIN trim_16
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  84.42 125.765 84.7 126.285 ;
    END
  END trim_16
  PIN trim_17
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  83.3 125.765 83.58 126.285 ;
    END
  END trim_17
  PIN trim_18
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  82.18 125.765 82.46 126.285 ;
    END
  END trim_18
  PIN trim_19
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  81.06 125.765 81.34 126.285 ;
    END
  END trim_19
  PIN trim_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  79.94 125.765 80.22 126.285 ;
    END
  END trim_2
  PIN trim_20
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  76.58 125.765 76.86 126.285 ;
    END
  END trim_20
  PIN trim_21
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  75.46 125.765 75.74 126.285 ;
    END
  END trim_21
  PIN trim_22
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  74.34 125.765 74.62 126.285 ;
    END
  END trim_22
  PIN trim_23
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  73.22 125.765 73.5 126.285 ;
    END
  END trim_23
  PIN trim_24
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  70.98 125.765 71.26 126.285 ;
    END
  END trim_24
  PIN trim_25
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  69.86 125.765 70.14 126.285 ;
    END
  END trim_25
  PIN trim_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  68.74 125.765 69.02 126.285 ;
    END
  END trim_3
  PIN trim_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  67.62 125.765 67.9 126.285 ;
    END
  END trim_4
  PIN trim_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  66.5 125.765 66.78 126.285 ;
    END
  END trim_5
  PIN trim_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  65.38 125.765 65.66 126.285 ;
    END
  END trim_6
  PIN trim_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  64.26 125.765 64.54 126.285 ;
    END
  END trim_7
  PIN trim_8
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  63.14 125.765 63.42 126.285 ;
    END
  END trim_8
  PIN trim_9
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  62.02 125.765 62.3 126.285 ;
    END
  END trim_9
  OBS
    LAYER Metal1 ;
     RECT  2.24 3.47 125.02 126.285 ;
    LAYER Metal2 ;
     RECT  2.24 3.47 125.02 126.285 ;
    LAYER Metal3 ;
     RECT  2.24 3.47 125.02 126.285 ;
    LAYER Metal4 ;
     RECT  2.24 3.47 125.02 126.285 ;
  END
END ring_osc2x13
END LIBRARY
