VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

VIA digital_pll_controller_via1_2_8960_1800_1_4_1240_1240
  VIARULE Via1_GEN_HH ;
  CUTSIZE 0.26 0.26 ;
  LAYERS Metal1 Via1 Metal2 ;
  CUTSPACING 0.36 0.36 ;
  ENCLOSURE 0.06 0.32 0.01 0.06 ;
  ROWCOL 1 4 ;
END digital_pll_controller_via1_2_8960_1800_1_4_1240_1240

VIA digital_pll_controller_via2_3_8960_560_1_8_1040_1040
  VIARULE Via2_GEN_HH ;
  CUTSIZE 0.26 0.26 ;
  LAYERS Metal2 Via2 Metal3 ;
  CUTSPACING 0.26 0.26 ;
  ENCLOSURE 0.01 0.06 0.06 0.01 ;
  ROWCOL 1 8 ;
END digital_pll_controller_via2_3_8960_560_1_8_1040_1040

VIA digital_pll_controller_via3_4_8960_560_1_8_1040_1040
  VIARULE Via3_GEN_HH ;
  CUTSIZE 0.26 0.26 ;
  LAYERS Metal3 Via3 Metal4 ;
  CUTSPACING 0.26 0.26 ;
  ENCLOSURE 0.06 0.01 0.29 0.06 ;
  ROWCOL 1 8 ;
END digital_pll_controller_via3_4_8960_560_1_8_1040_1040

MACRO digital_pll_controller
  FOREIGN digital_pll_controller 0 0 ;
  CLASS BLOCK ;
  SIZE 162.805 BY 162.805 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER Metal4 ;
        RECT  117.04 7.39 121.52 157.25 ;
        RECT  72.24 7.39 76.72 157.25 ;
        RECT  27.44 7.39 31.92 157.25 ;
      LAYER Metal1 ;
        RECT  2.24 156.35 160.72 157.25 ;
        RECT  2.24 148.51 160.72 149.41 ;
        RECT  2.24 140.67 160.72 141.57 ;
        RECT  2.24 132.83 160.72 133.73 ;
        RECT  2.24 124.99 160.72 125.89 ;
        RECT  2.24 117.15 160.72 118.05 ;
        RECT  2.24 109.31 160.72 110.21 ;
        RECT  2.24 101.47 160.72 102.37 ;
        RECT  2.24 93.63 160.72 94.53 ;
        RECT  2.24 85.79 160.72 86.69 ;
        RECT  2.24 77.95 160.72 78.85 ;
        RECT  2.24 70.11 160.72 71.01 ;
        RECT  2.24 62.27 160.72 63.17 ;
        RECT  2.24 54.43 160.72 55.33 ;
        RECT  2.24 46.59 160.72 47.49 ;
        RECT  2.24 38.75 160.72 39.65 ;
        RECT  2.24 30.91 160.72 31.81 ;
        RECT  2.24 23.07 160.72 23.97 ;
        RECT  2.24 15.23 160.72 16.13 ;
        RECT  2.24 7.39 160.72 8.29 ;
      VIA 119.28 156.8 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 156.8 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 156.8 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 148.96 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 148.96 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 148.96 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 141.12 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 141.12 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 141.12 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 133.28 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 133.28 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 133.28 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 125.44 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 125.44 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 125.44 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 117.6 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 117.6 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 117.6 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 109.76 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 109.76 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 109.76 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 101.92 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 101.92 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 101.92 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 94.08 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 94.08 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 94.08 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 86.24 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 86.24 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 86.24 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 78.4 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 78.4 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 78.4 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 70.56 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 70.56 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 70.56 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 62.72 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 62.72 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 62.72 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 54.88 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 54.88 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 54.88 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 47.04 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 47.04 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 47.04 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 39.2 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 39.2 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 39.2 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 31.36 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 31.36 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 31.36 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 23.52 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 23.52 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 23.52 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 15.68 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 15.68 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 15.68 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 7.84 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 7.84 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 7.84 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 156.8 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 156.8 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 156.8 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 148.96 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 148.96 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 148.96 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 141.12 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 141.12 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 141.12 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 133.28 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 133.28 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 133.28 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 125.44 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 125.44 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 125.44 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 117.6 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 117.6 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 117.6 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 109.76 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 109.76 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 109.76 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 101.92 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 101.92 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 101.92 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 94.08 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 94.08 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 94.08 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 86.24 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 86.24 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 86.24 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 78.4 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 78.4 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 78.4 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 70.56 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 70.56 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 70.56 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 62.72 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 62.72 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 62.72 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 54.88 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 54.88 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 54.88 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 47.04 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 47.04 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 47.04 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 39.2 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 39.2 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 39.2 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 31.36 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 31.36 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 31.36 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 23.52 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 23.52 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 23.52 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 15.68 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 15.68 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 15.68 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 7.84 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 7.84 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 7.84 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 156.8 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 156.8 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 156.8 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 148.96 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 148.96 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 148.96 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 141.12 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 141.12 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 141.12 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 133.28 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 133.28 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 133.28 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 125.44 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 125.44 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 125.44 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 117.6 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 117.6 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 117.6 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 109.76 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 109.76 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 109.76 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 101.92 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 101.92 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 101.92 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 94.08 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 94.08 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 94.08 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 86.24 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 86.24 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 86.24 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 78.4 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 78.4 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 78.4 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 70.56 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 70.56 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 70.56 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 62.72 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 62.72 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 62.72 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 54.88 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 54.88 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 54.88 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 47.04 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 47.04 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 47.04 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 39.2 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 39.2 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 39.2 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 31.36 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 31.36 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 31.36 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 23.52 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 23.52 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 23.52 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 15.68 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 15.68 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 15.68 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 7.84 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 7.84 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 7.84 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER Metal4 ;
        RECT  156.8 3.47 161.28 161.17 ;
        RECT  112 3.47 116.48 161.17 ;
        RECT  67.2 3.47 71.68 161.17 ;
        RECT  22.4 3.47 26.88 161.17 ;
      LAYER Metal1 ;
        RECT  2.24 160.27 161.28 161.17 ;
        RECT  2.24 152.43 161.28 153.33 ;
        RECT  2.24 144.59 161.28 145.49 ;
        RECT  2.24 136.75 161.28 137.65 ;
        RECT  2.24 128.91 161.28 129.81 ;
        RECT  2.24 121.07 161.28 121.97 ;
        RECT  2.24 113.23 161.28 114.13 ;
        RECT  2.24 105.39 161.28 106.29 ;
        RECT  2.24 97.55 161.28 98.45 ;
        RECT  2.24 89.71 161.28 90.61 ;
        RECT  2.24 81.87 161.28 82.77 ;
        RECT  2.24 74.03 161.28 74.93 ;
        RECT  2.24 66.19 161.28 67.09 ;
        RECT  2.24 58.35 161.28 59.25 ;
        RECT  2.24 50.51 161.28 51.41 ;
        RECT  2.24 42.67 161.28 43.57 ;
        RECT  2.24 34.83 161.28 35.73 ;
        RECT  2.24 26.99 161.28 27.89 ;
        RECT  2.24 19.15 161.28 20.05 ;
        RECT  2.24 11.31 161.28 12.21 ;
        RECT  2.24 3.47 161.28 4.37 ;
      VIA 159.04 160.72 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 160.72 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 160.72 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 152.88 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 152.88 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 152.88 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 145.04 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 145.04 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 145.04 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 137.2 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 137.2 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 137.2 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 129.36 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 129.36 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 129.36 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 121.52 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 121.52 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 121.52 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 113.68 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 113.68 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 113.68 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 105.84 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 105.84 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 105.84 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 98 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 98 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 98 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 90.16 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 90.16 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 90.16 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 82.32 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 82.32 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 82.32 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 74.48 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 74.48 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 74.48 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 66.64 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 66.64 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 66.64 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 58.8 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 58.8 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 58.8 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 50.96 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 50.96 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 50.96 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 43.12 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 43.12 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 43.12 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 35.28 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 35.28 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 35.28 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 27.44 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 27.44 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 27.44 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 19.6 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 19.6 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 19.6 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 11.76 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 11.76 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 11.76 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 159.04 3.92 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 159.04 3.92 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 159.04 3.92 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 160.72 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 160.72 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 160.72 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 152.88 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 152.88 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 152.88 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 145.04 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 145.04 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 145.04 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 137.2 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 137.2 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 137.2 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 129.36 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 129.36 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 129.36 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 121.52 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 121.52 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 121.52 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 113.68 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 113.68 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 113.68 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 105.84 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 105.84 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 105.84 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 98 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 98 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 98 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 90.16 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 90.16 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 90.16 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 82.32 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 82.32 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 82.32 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 74.48 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 74.48 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 74.48 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 66.64 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 66.64 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 66.64 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 58.8 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 58.8 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 58.8 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 50.96 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 50.96 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 50.96 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 43.12 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 43.12 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 43.12 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 35.28 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 35.28 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 35.28 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 27.44 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 27.44 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 27.44 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 19.6 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 19.6 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 19.6 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 11.76 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 11.76 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 11.76 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 3.92 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 3.92 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 3.92 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 160.72 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 160.72 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 160.72 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 152.88 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 152.88 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 152.88 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 145.04 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 145.04 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 145.04 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 137.2 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 137.2 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 137.2 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 129.36 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 129.36 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 129.36 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 121.52 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 121.52 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 121.52 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 113.68 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 113.68 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 113.68 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 105.84 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 105.84 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 105.84 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 98 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 98 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 98 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 90.16 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 90.16 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 90.16 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 82.32 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 82.32 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 82.32 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 74.48 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 74.48 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 74.48 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 66.64 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 66.64 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 66.64 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 58.8 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 58.8 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 58.8 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 50.96 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 50.96 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 50.96 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 43.12 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 43.12 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 43.12 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 35.28 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 35.28 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 35.28 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 27.44 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 27.44 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 27.44 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 19.6 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 19.6 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 19.6 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 11.76 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 11.76 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 11.76 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 3.92 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 3.92 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 3.92 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 160.72 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 160.72 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 160.72 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 152.88 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 152.88 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 152.88 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 145.04 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 145.04 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 145.04 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 137.2 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 137.2 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 137.2 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 129.36 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 129.36 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 129.36 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 121.52 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 121.52 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 121.52 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 113.68 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 113.68 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 113.68 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 105.84 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 105.84 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 105.84 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 98 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 98 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 98 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 90.16 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 90.16 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 90.16 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 82.32 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 82.32 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 82.32 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 74.48 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 74.48 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 74.48 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 66.64 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 66.64 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 66.64 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 58.8 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 58.8 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 58.8 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 50.96 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 50.96 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 50.96 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 43.12 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 43.12 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 43.12 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 35.28 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 35.28 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 35.28 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 27.44 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 27.44 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 27.44 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 19.6 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 19.6 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 19.6 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 11.76 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 11.76 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 11.76 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 3.92 digital_pll_controller_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 3.92 digital_pll_controller_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 3.92 digital_pll_controller_via1_2_8960_1800_1_4_1240_1240 ;
    END
  END VSS
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  100.1 162.285 100.38 162.805 ;
    END
  END clock
  PIN dco
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  29.54 162.285 29.82 162.805 ;
    END
  END dco
  PIN div[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  87.78 162.285 88.06 162.805 ;
    END
  END div[0]
  PIN div[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  83.3 162.285 83.58 162.805 ;
    END
  END div[1]
  PIN div[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  90.02 162.285 90.3 162.805 ;
    END
  END div[2]
  PIN div[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  88.9 162.285 89.18 162.805 ;
    END
  END div[3]
  PIN div[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  91.14 162.285 91.42 162.805 ;
    END
  END div[4]
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  27.3 162.285 27.58 162.805 ;
    END
  END enable
  PIN osc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  11.62 162.285 11.9 162.805 ;
    END
  END osc
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  28.42 162.285 28.7 162.805 ;
    END
  END reset
  PIN trim[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  119.14 162.285 119.42 162.805 ;
    END
  END trim[0]
  PIN trim[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  124.74 162.285 125.02 162.805 ;
    END
  END trim[10]
  PIN trim[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  142.66 162.285 142.94 162.805 ;
    END
  END trim[11]
  PIN trim[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  128.1 162.285 128.38 162.805 ;
    END
  END trim[12]
  PIN trim[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  140.42 162.285 140.7 162.805 ;
    END
  END trim[13]
  PIN trim[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  113.54 162.285 113.82 162.805 ;
    END
  END trim[14]
  PIN trim[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  139.3 162.285 139.58 162.805 ;
    END
  END trim[15]
  PIN trim[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  125.86 162.285 126.14 162.805 ;
    END
  END trim[16]
  PIN trim[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  141.54 162.285 141.82 162.805 ;
    END
  END trim[17]
  PIN trim[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  126.98 162.285 127.26 162.805 ;
    END
  END trim[18]
  PIN trim[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  137.06 162.285 137.34 162.805 ;
    END
  END trim[19]
  PIN trim[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  132.58 162.285 132.86 162.805 ;
    END
  END trim[1]
  PIN trim[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  110.18 162.285 110.46 162.805 ;
    END
  END trim[20]
  PIN trim[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  133.7 162.285 133.98 162.805 ;
    END
  END trim[21]
  PIN trim[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  138.18 162.285 138.46 162.805 ;
    END
  END trim[22]
  PIN trim[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  129.22 162.285 129.5 162.805 ;
    END
  END trim[23]
  PIN trim[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  111.3 162.285 111.58 162.805 ;
    END
  END trim[24]
  PIN trim[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  135.94 162.285 136.22 162.805 ;
    END
  END trim[25]
  PIN trim[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  121.38 162.285 121.66 162.805 ;
    END
  END trim[2]
  PIN trim[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  122.5 162.285 122.78 162.805 ;
    END
  END trim[3]
  PIN trim[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  112.42 162.285 112.7 162.805 ;
    END
  END trim[4]
  PIN trim[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  130.34 162.285 130.62 162.805 ;
    END
  END trim[5]
  PIN trim[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  123.62 162.285 123.9 162.805 ;
    END
  END trim[6]
  PIN trim[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  134.82 162.285 135.1 162.805 ;
    END
  END trim[7]
  PIN trim[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  131.46 162.285 131.74 162.805 ;
    END
  END trim[8]
  PIN trim[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  115.78 162.285 116.06 162.805 ;
    END
  END trim[9]
  OBS
    LAYER Metal1 ;
     RECT  2.24 3.47 161.28 162.805 ;
    LAYER Metal2 ;
     RECT  2.24 3.47 161.28 162.805 ;
    LAYER Metal3 ;
     RECT  2.24 3.47 161.28 162.805 ;
    LAYER Metal4 ;
     RECT  2.24 3.47 161.28 162.805 ;
  END
END digital_pll_controller
END LIBRARY
