module digital_pll (dco,
    enable,
    osc,
    resetb,
    clockp,
    div,
    ext_trim);
 input dco;
 input enable;
 input osc;
 input resetb;
 output [1:0] clockp;
 input [4:0] div;
 input [25:0] ext_trim;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire net33;
 wire net32;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire net31;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire net30;
 wire _168_;
 wire net29;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire net28;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire net35;
 wire net36;
 wire ireset;
 wire \itrim[0] ;
 wire \itrim[10] ;
 wire \itrim[11] ;
 wire \itrim[12] ;
 wire \itrim[13] ;
 wire \itrim[14] ;
 wire \itrim[15] ;
 wire \itrim[16] ;
 wire \itrim[17] ;
 wire \itrim[18] ;
 wire \itrim[19] ;
 wire \itrim[1] ;
 wire \itrim[20] ;
 wire \itrim[21] ;
 wire \itrim[22] ;
 wire \itrim[23] ;
 wire \itrim[24] ;
 wire \itrim[25] ;
 wire \itrim[2] ;
 wire \itrim[3] ;
 wire \itrim[4] ;
 wire \itrim[5] ;
 wire \itrim[6] ;
 wire \itrim[7] ;
 wire \itrim[8] ;
 wire \itrim[9] ;
 wire net27;
 wire \pll_control.count0[0] ;
 wire \pll_control.count0[1] ;
 wire \pll_control.count0[2] ;
 wire \pll_control.count0[3] ;
 wire \pll_control.count0[4] ;
 wire \pll_control.count1[0] ;
 wire \pll_control.count1[1] ;
 wire \pll_control.count1[2] ;
 wire \pll_control.count1[3] ;
 wire \pll_control.count1[4] ;
 wire \pll_control.oscbuf[0] ;
 wire \pll_control.oscbuf[1] ;
 wire \pll_control.oscbuf[2] ;
 wire \pll_control.prep[0] ;
 wire \pll_control.prep[1] ;
 wire \pll_control.prep[2] ;
 wire \pll_control.tint[0] ;
 wire \pll_control.tint[1] ;
 wire \pll_control.tint[2] ;
 wire \pll_control.tint[3] ;
 wire \pll_control.tint[4] ;
 wire \pll_control.tval[0] ;
 wire \pll_control.tval[1] ;
 wire \ringosc.c[0] ;
 wire \ringosc.c[1] ;
 wire net25;
 wire \ringosc.dstage[0].id.d1 ;
 wire \ringosc.dstage[0].id.d2 ;
 wire \ringosc.dstage[0].id.in ;
 wire \ringosc.dstage[0].id.out ;
 wire \ringosc.dstage[0].id.trim0b ;
 wire \ringosc.dstage[0].id.trim1b ;
 wire net26;
 wire net23;
 wire \ringosc.dstage[10].id.d1 ;
 wire \ringosc.dstage[10].id.d2 ;
 wire \ringosc.dstage[10].id.in ;
 wire \ringosc.dstage[10].id.out ;
 wire \ringosc.dstage[10].id.trim0b ;
 wire \ringosc.dstage[10].id.trim1b ;
 wire net24;
 wire net21;
 wire \ringosc.dstage[11].id.d1 ;
 wire \ringosc.dstage[11].id.d2 ;
 wire \ringosc.dstage[11].id.out ;
 wire \ringosc.dstage[11].id.trim0b ;
 wire \ringosc.dstage[11].id.trim1b ;
 wire net22;
 wire net19;
 wire \ringosc.dstage[1].id.d1 ;
 wire \ringosc.dstage[1].id.d2 ;
 wire \ringosc.dstage[1].id.out ;
 wire \ringosc.dstage[1].id.trim0b ;
 wire \ringosc.dstage[1].id.trim1b ;
 wire net20;
 wire net17;
 wire \ringosc.dstage[2].id.d1 ;
 wire \ringosc.dstage[2].id.d2 ;
 wire \ringosc.dstage[2].id.out ;
 wire \ringosc.dstage[2].id.trim0b ;
 wire \ringosc.dstage[2].id.trim1b ;
 wire net18;
 wire net15;
 wire \ringosc.dstage[3].id.d1 ;
 wire \ringosc.dstage[3].id.d2 ;
 wire \ringosc.dstage[3].id.out ;
 wire \ringosc.dstage[3].id.trim0b ;
 wire \ringosc.dstage[3].id.trim1b ;
 wire net16;
 wire net13;
 wire \ringosc.dstage[4].id.d1 ;
 wire \ringosc.dstage[4].id.d2 ;
 wire \ringosc.dstage[4].id.out ;
 wire \ringosc.dstage[4].id.trim0b ;
 wire \ringosc.dstage[4].id.trim1b ;
 wire net14;
 wire net11;
 wire \ringosc.dstage[5].id.d1 ;
 wire \ringosc.dstage[5].id.d2 ;
 wire \ringosc.dstage[5].id.out ;
 wire \ringosc.dstage[5].id.trim0b ;
 wire \ringosc.dstage[5].id.trim1b ;
 wire net12;
 wire net9;
 wire \ringosc.dstage[6].id.d1 ;
 wire \ringosc.dstage[6].id.d2 ;
 wire \ringosc.dstage[6].id.out ;
 wire \ringosc.dstage[6].id.trim0b ;
 wire \ringosc.dstage[6].id.trim1b ;
 wire net10;
 wire net7;
 wire \ringosc.dstage[7].id.d1 ;
 wire \ringosc.dstage[7].id.d2 ;
 wire \ringosc.dstage[7].id.out ;
 wire \ringosc.dstage[7].id.trim0b ;
 wire \ringosc.dstage[7].id.trim1b ;
 wire net8;
 wire net5;
 wire \ringosc.dstage[8].id.d1 ;
 wire \ringosc.dstage[8].id.d2 ;
 wire \ringosc.dstage[8].id.out ;
 wire \ringosc.dstage[8].id.trim0b ;
 wire \ringosc.dstage[8].id.trim1b ;
 wire net6;
 wire net3;
 wire \ringosc.dstage[9].id.d1 ;
 wire \ringosc.dstage[9].id.d2 ;
 wire \ringosc.dstage[9].id.trim0b ;
 wire \ringosc.dstage[9].id.trim1b ;
 wire net4;
 wire \ringosc.iss.ctrl0b ;
 wire net2;
 wire \ringosc.iss.d1 ;
 wire \ringosc.iss.d2 ;
 wire \ringosc.iss.trim1b ;
 wire net1;
 wire net34;

 gf180mcu_fd_sc_mcu7t5v0__and3_2 _278_ (.A1(\pll_control.count0[2] ),
    .A2(\pll_control.count0[3] ),
    .A3(_032_),
    .Z(_034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _279_ (.A1(net7),
    .A2(net34),
    .ZN(ireset));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input32 (.I(ext_trim[9]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input31 (.I(ext_trim[8]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _282_ (.A1(ireset),
    .A2(net2),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _283_ (.I(net6),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _284_ (.A1(_001_),
    .A2(_008_),
    .A3(_010_),
    .Z(_070_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _285_ (.A1(_008_),
    .A2(_009_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _286_ (.A1(_070_),
    .A2(_007_),
    .A3(_071_),
    .Z(_072_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _287_ (.A1(_006_),
    .A2(_072_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _288_ (.I(net5),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _289_ (.I(net4),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _290_ (.I(net3),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _291_ (.A1(_023_),
    .A2(_020_),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _292_ (.I(_019_),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _293_ (.A1(_073_),
    .A2(_074_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _294_ (.A1(_075_),
    .A2(_016_),
    .B(_015_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _295_ (.I(_030_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _296_ (.A1(_077_),
    .A2(_027_),
    .B(_026_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _297_ (.A1(_016_),
    .A2(_020_),
    .A3(_024_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _298_ (.A1(_078_),
    .A2(_079_),
    .Z(_080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _299_ (.A1(_076_),
    .A2(_080_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _300_ (.A1(_027_),
    .A2(_031_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _301_ (.A1(_079_),
    .A2(_082_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _302_ (.I(_083_),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _303_ (.A1(_081_),
    .A2(_084_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _304_ (.A1(_010_),
    .A2(_011_),
    .B(_009_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _305_ (.A1(_000_),
    .A2(_010_),
    .A3(_012_),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _306_ (.A1(_086_),
    .A2(_087_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _307_ (.A1(_006_),
    .A2(_008_),
    .Z(_089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _308_ (.A1(_088_),
    .A2(_089_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _309_ (.A1(_006_),
    .A2(_007_),
    .B(_005_),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _310_ (.A1(_090_),
    .A2(_091_),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _311_ (.I(_092_),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _312_ (.A1(_085_),
    .A2(_093_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _313_ (.A1(_008_),
    .A2(_088_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _314_ (.A1(_001_),
    .A2(_010_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _315_ (.I(_028_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _316_ (.I(_035_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _317_ (.A1(\pll_control.count0[0] ),
    .A2(_094_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _318_ (.I(\pll_control.oscbuf[1] ),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _319_ (.A1(_096_),
    .A2(\pll_control.oscbuf[2] ),
    .Z(_097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _320_ (.A1(_096_),
    .A2(\pll_control.oscbuf[2] ),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _321_ (.A1(_097_),
    .A2(_098_),
    .Z(_099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input30 (.I(ext_trim[7]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _323_ (.A1(_095_),
    .A2(_099_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _324_ (.I0(_033_),
    .I1(\pll_control.count0[1] ),
    .S(_035_),
    .Z(_101_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _325_ (.A1(_101_),
    .A2(_099_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _326_ (.I(_032_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _327_ (.I(\pll_control.count0[2] ),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _328_ (.A1(_102_),
    .A2(_035_),
    .B(_103_),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _329_ (.A1(_103_),
    .A2(_102_),
    .A3(_035_),
    .Z(_105_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _330_ (.A1(_099_),
    .A2(_104_),
    .A3(_105_),
    .Z(_050_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _331_ (.A1(_094_),
    .A2(\pll_control.count0[2] ),
    .A3(\pll_control.count0[0] ),
    .A4(\pll_control.count0[1] ),
    .Z(_106_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _332_ (.A1(_106_),
    .A2(\pll_control.count0[3] ),
    .Z(_107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _333_ (.A1(_106_),
    .A2(\pll_control.count0[3] ),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _334_ (.A1(_107_),
    .A2(_099_),
    .A3(_108_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _335_ (.I0(_036_),
    .I1(\pll_control.count0[4] ),
    .S(_035_),
    .Z(_109_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _336_ (.A1(_109_),
    .A2(_099_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _337_ (.A1(\pll_control.tint[3] ),
    .A2(\pll_control.tint[4] ),
    .Z(_110_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _338_ (.A1(_110_),
    .A2(\pll_control.tval[0] ),
    .A3(\pll_control.tval[1] ),
    .Z(_111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _339_ (.A1(\pll_control.tint[1] ),
    .A2(\pll_control.tint[0] ),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _340_ (.I(_112_),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _341_ (.A1(_111_),
    .A2(\pll_control.tint[2] ),
    .A3(_113_),
    .ZN(_114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _342_ (.A1(_002_),
    .A2(_114_),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _343_ (.I(_115_),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _344_ (.I(_099_),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu7t5v0__and4_4 _345_ (.A1(_117_),
    .A2(\pll_control.prep[1] ),
    .A3(\pll_control.prep[0] ),
    .A4(\pll_control.prep[2] ),
    .Z(_118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _346_ (.I(_081_),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _347_ (.I(\pll_control.tint[3] ),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _348_ (.I(\pll_control.tint[2] ),
    .ZN(_121_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _349_ (.A1(_120_),
    .A2(_121_),
    .Z(_122_));
 gf180mcu_fd_sc_mcu7t5v0__inv_8 _350_ (.I(\pll_control.tint[4] ),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _351_ (.A1(_122_),
    .A2(_123_),
    .ZN(_124_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _352_ (.A1(\pll_control.tval[0] ),
    .A2(\pll_control.tval[1] ),
    .Z(_125_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _353_ (.I(\pll_control.tint[1] ),
    .ZN(_126_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _354_ (.I(\pll_control.tint[0] ),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _355_ (.A1(_126_),
    .A2(_127_),
    .Z(_128_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _356_ (.I(_128_),
    .ZN(_129_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _357_ (.A1(_124_),
    .A2(_125_),
    .A3(_129_),
    .Z(_130_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _358_ (.A1(_093_),
    .A2(_119_),
    .A3(_130_),
    .ZN(_131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _359_ (.A1(_002_),
    .A2(_131_),
    .ZN(_132_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _360_ (.A1(_116_),
    .A2(_118_),
    .A3(_132_),
    .ZN(_133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _361_ (.A1(_133_),
    .A2(\pll_control.tval[0] ),
    .ZN(_134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _362_ (.A1(_132_),
    .A2(_118_),
    .ZN(_135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _363_ (.A1(_135_),
    .A2(_115_),
    .ZN(_136_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _364_ (.I(\pll_control.tval[0] ),
    .ZN(_137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _365_ (.A1(_136_),
    .A2(_137_),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _366_ (.A1(_134_),
    .A2(_138_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _367_ (.A1(_133_),
    .A2(\pll_control.tval[1] ),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _368_ (.A1(_136_),
    .A2(_004_),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _369_ (.A1(_139_),
    .A2(_140_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _370_ (.A1(_133_),
    .A2(\pll_control.tint[0] ),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _371_ (.I(_040_),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _372_ (.A1(_003_),
    .A2(_142_),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _373_ (.A1(_136_),
    .A2(_143_),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _374_ (.A1(_141_),
    .A2(_144_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _375_ (.A1(_133_),
    .A2(\pll_control.tint[1] ),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _376_ (.I(_042_),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _377_ (.I(_038_),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _378_ (.A1(_040_),
    .A2(_037_),
    .B(_039_),
    .ZN(_148_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _379_ (.A1(_137_),
    .A2(_147_),
    .A3(_142_),
    .B(_148_),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _380_ (.A1(_146_),
    .A2(_149_),
    .ZN(_150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _381_ (.A1(_136_),
    .A2(_150_),
    .ZN(_151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _382_ (.A1(_145_),
    .A2(_151_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _383_ (.A1(_133_),
    .A2(\pll_control.tint[2] ),
    .ZN(_152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _384_ (.I(_044_),
    .ZN(_153_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _385_ (.I(_003_),
    .ZN(_154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _386_ (.A1(_042_),
    .A2(_039_),
    .B(_041_),
    .ZN(_155_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _387_ (.A1(_154_),
    .A2(_142_),
    .A3(_146_),
    .B(_155_),
    .ZN(_156_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _388_ (.A1(_153_),
    .A2(_156_),
    .ZN(_157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _389_ (.A1(_136_),
    .A2(_157_),
    .ZN(_158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _390_ (.A1(_152_),
    .A2(_158_),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _391_ (.A1(_133_),
    .A2(\pll_control.tint[3] ),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _392_ (.A1(_042_),
    .A2(_044_),
    .ZN(_160_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _393_ (.A1(_160_),
    .A2(_137_),
    .A3(_147_),
    .A4(_142_),
    .Z(_161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _394_ (.A1(_044_),
    .A2(_041_),
    .B(_043_),
    .ZN(_162_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _395_ (.A1(_148_),
    .A2(_160_),
    .B(_161_),
    .C(_162_),
    .ZN(_163_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _396_ (.A1(_046_),
    .A2(_163_),
    .Z(_164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _397_ (.A1(_136_),
    .A2(_164_),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _398_ (.A1(_159_),
    .A2(_165_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _399_ (.A1(_076_),
    .A2(_080_),
    .B(_083_),
    .ZN(_166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input29 (.I(ext_trim[6]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _401_ (.A1(_166_),
    .A2(_092_),
    .B(_123_),
    .ZN(_168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input28 (.I(ext_trim[5]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _403_ (.A1(_085_),
    .A2(\pll_control.tint[4] ),
    .A3(_093_),
    .ZN(_170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _404_ (.A1(_168_),
    .A2(_170_),
    .ZN(_171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _405_ (.A1(_044_),
    .A2(_046_),
    .ZN(_172_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _406_ (.A1(_172_),
    .A2(_154_),
    .A3(_142_),
    .A4(_146_),
    .Z(_173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _407_ (.A1(_046_),
    .A2(_043_),
    .B(_045_),
    .ZN(_174_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _408_ (.A1(_155_),
    .A2(_172_),
    .Z(_175_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _409_ (.A1(_173_),
    .A2(_174_),
    .A3(_175_),
    .Z(_176_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _410_ (.I(_176_),
    .ZN(_177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _411_ (.A1(_171_),
    .A2(_177_),
    .ZN(_178_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _412_ (.A1(_168_),
    .A2(_170_),
    .A3(_176_),
    .ZN(_179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _413_ (.A1(_178_),
    .A2(_179_),
    .ZN(_180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _414_ (.A1(_180_),
    .A2(_136_),
    .ZN(_181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _415_ (.A1(_133_),
    .A2(\pll_control.tint[4] ),
    .ZN(_182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _416_ (.A1(_181_),
    .A2(_182_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _417_ (.I0(\pll_control.count0[0] ),
    .I1(\pll_control.count1[0] ),
    .S(_099_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _418_ (.I0(\pll_control.count0[1] ),
    .I1(\pll_control.count1[1] ),
    .S(_099_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _419_ (.I0(\pll_control.count0[2] ),
    .I1(\pll_control.count1[2] ),
    .S(_099_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _420_ (.I0(\pll_control.count0[3] ),
    .I1(\pll_control.count1[3] ),
    .S(_099_),
    .Z(_056_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _421_ (.I0(\pll_control.count0[4] ),
    .I1(\pll_control.count1[4] ),
    .S(_099_),
    .Z(_057_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _422_ (.A1(_117_),
    .A2(\pll_control.prep[0] ),
    .Z(_058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _423_ (.I0(\pll_control.prep[0] ),
    .I1(\pll_control.prep[1] ),
    .S(_099_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _424_ (.I0(\pll_control.prep[1] ),
    .I1(\pll_control.prep[2] ),
    .S(_099_),
    .Z(_060_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _425_ (.A1(_122_),
    .A2(_128_),
    .Z(_183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _426_ (.A1(_183_),
    .A2(_123_),
    .ZN(_184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _427_ (.I0(_184_),
    .I1(net8),
    .S(net2),
    .Z(\itrim[0] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _428_ (.I(net2),
    .ZN(_185_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _429_ (.A1(_124_),
    .A2(_185_),
    .Z(_186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _430_ (.A1(_185_),
    .A2(_113_),
    .B(_186_),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _431_ (.A1(net2),
    .A2(net9),
    .ZN(_188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _432_ (.A1(_187_),
    .A2(_188_),
    .ZN(\itrim[10] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _433_ (.A1(_120_),
    .A2(\pll_control.tint[2] ),
    .Z(_189_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _434_ (.A1(_189_),
    .A2(_113_),
    .Z(_190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _435_ (.A1(_190_),
    .A2(_123_),
    .ZN(_191_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _436_ (.A1(_128_),
    .A2(_189_),
    .Z(_192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _437_ (.A1(_192_),
    .A2(_123_),
    .ZN(_193_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _438_ (.A1(_186_),
    .A2(_193_),
    .Z(_194_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _439_ (.A1(_123_),
    .A2(_127_),
    .A3(\pll_control.tint[1] ),
    .Z(_195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _440_ (.A1(_126_),
    .A2(\pll_control.tint[0] ),
    .ZN(_196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _441_ (.A1(_196_),
    .A2(\pll_control.tint[4] ),
    .ZN(_197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _442_ (.A1(_195_),
    .A2(_197_),
    .B(_189_),
    .ZN(_198_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _443_ (.A1(_194_),
    .A2(_198_),
    .Z(_199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _444_ (.A1(_121_),
    .A2(\pll_control.tint[3] ),
    .ZN(_200_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _445_ (.A1(_196_),
    .A2(_200_),
    .A3(\pll_control.tint[4] ),
    .Z(_201_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _446_ (.A1(_129_),
    .A2(_200_),
    .A3(\pll_control.tint[4] ),
    .Z(_202_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _447_ (.A1(_191_),
    .A2(_199_),
    .A3(_201_),
    .A4(_202_),
    .ZN(_203_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _448_ (.I(_200_),
    .ZN(_204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _449_ (.A1(_195_),
    .A2(_204_),
    .ZN(_205_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _450_ (.I(_205_),
    .ZN(_206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input27 (.I(ext_trim[4]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _452_ (.A1(net2),
    .A2(net10),
    .ZN(_208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _453_ (.A1(_203_),
    .A2(_206_),
    .B(_208_),
    .ZN(\itrim[11] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _454_ (.I(_194_),
    .ZN(_209_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _455_ (.A1(_197_),
    .A2(_189_),
    .Z(_210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _456_ (.A1(net2),
    .A2(net11),
    .ZN(_211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _457_ (.A1(_209_),
    .A2(_210_),
    .B(_211_),
    .ZN(\itrim[12] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _458_ (.A1(_202_),
    .A2(_191_),
    .Z(_212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _459_ (.A1(_199_),
    .A2(_212_),
    .ZN(_213_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _460_ (.I(_213_),
    .ZN(_214_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _461_ (.A1(\pll_control.tint[3] ),
    .A2(\pll_control.tint[2] ),
    .Z(_215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _462_ (.A1(\pll_control.tint[0] ),
    .A2(_204_),
    .B1(_128_),
    .B2(_215_),
    .ZN(_216_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _463_ (.A1(_216_),
    .A2(\pll_control.tint[4] ),
    .ZN(_217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _464_ (.A1(_217_),
    .A2(_206_),
    .ZN(_218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _465_ (.A1(_214_),
    .A2(_218_),
    .ZN(_219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _466_ (.A1(_197_),
    .A2(_215_),
    .ZN(_220_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _467_ (.I(_220_),
    .ZN(_221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _468_ (.A1(net2),
    .A2(net12),
    .ZN(_222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _469_ (.A1(_219_),
    .A2(_221_),
    .B(_222_),
    .ZN(\itrim[13] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _470_ (.A1(_122_),
    .A2(\pll_control.tint[4] ),
    .Z(_223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _471_ (.A1(_223_),
    .A2(_112_),
    .ZN(_224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _472_ (.A1(_113_),
    .A2(_215_),
    .ZN(_225_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _473_ (.A1(_225_),
    .A2(\pll_control.tint[4] ),
    .Z(_226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _474_ (.A1(_195_),
    .A2(_215_),
    .ZN(_227_));
 gf180mcu_fd_sc_mcu7t5v0__and4_4 _475_ (.A1(_224_),
    .A2(_220_),
    .A3(_226_),
    .A4(_227_),
    .Z(_228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _476_ (.A1(_228_),
    .A2(_218_),
    .ZN(_229_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _477_ (.I(_189_),
    .ZN(_230_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _478_ (.A1(_122_),
    .A2(_113_),
    .Z(_231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _479_ (.A1(_231_),
    .A2(\pll_control.tint[4] ),
    .ZN(_232_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _480_ (.A1(_123_),
    .A2(\pll_control.tint[1] ),
    .A3(_230_),
    .B(_232_),
    .ZN(_233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _481_ (.A1(_229_),
    .A2(_233_),
    .ZN(_234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _482_ (.A1(_234_),
    .A2(_199_),
    .ZN(_235_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _483_ (.A1(_230_),
    .A2(_123_),
    .A3(_126_),
    .A4(\pll_control.tint[0] ),
    .Z(_236_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _484_ (.I(_190_),
    .ZN(_237_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _485_ (.A1(_129_),
    .A2(_200_),
    .B(_236_),
    .C(_237_),
    .ZN(_238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _486_ (.A1(net2),
    .A2(net13),
    .ZN(_239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _487_ (.A1(_235_),
    .A2(_238_),
    .B(_239_),
    .ZN(\itrim[14] ));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _488_ (.A1(_198_),
    .A2(_228_),
    .A3(_218_),
    .A4(_212_),
    .ZN(_240_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _489_ (.A1(_129_),
    .A2(_230_),
    .B(_186_),
    .C(_232_),
    .ZN(_241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _490_ (.A1(net2),
    .A2(net14),
    .ZN(_242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _491_ (.A1(_240_),
    .A2(_241_),
    .B(_242_),
    .ZN(\itrim[15] ));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _492_ (.A1(_183_),
    .A2(_123_),
    .A3(net2),
    .Z(_243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _493_ (.A1(net2),
    .A2(net15),
    .ZN(_244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _494_ (.A1(_243_),
    .A2(_244_),
    .ZN(\itrim[16] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _495_ (.A1(_234_),
    .A2(_214_),
    .A3(_236_),
    .ZN(_245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _496_ (.A1(net2),
    .A2(net16),
    .ZN(_246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _497_ (.A1(_245_),
    .A2(_246_),
    .ZN(\itrim[17] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _498_ (.I(_193_),
    .ZN(_247_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _499_ (.A1(_187_),
    .A2(_231_),
    .A3(_247_),
    .Z(_248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _500_ (.A1(net2),
    .A2(net17),
    .ZN(_249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _501_ (.A1(_240_),
    .A2(_248_),
    .B(_249_),
    .ZN(\itrim[18] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _502_ (.A1(_225_),
    .A2(_123_),
    .ZN(_250_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _503_ (.I0(_250_),
    .I1(net18),
    .S(net2),
    .Z(\itrim[19] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _504_ (.I(_199_),
    .ZN(_251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _505_ (.A1(_237_),
    .A2(_200_),
    .B(\pll_control.tint[4] ),
    .ZN(_252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _506_ (.A1(net2),
    .A2(net19),
    .ZN(_253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _507_ (.A1(_251_),
    .A2(_252_),
    .B(_253_),
    .ZN(\itrim[1] ));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _508_ (.A1(\pll_control.tint[1] ),
    .A2(\pll_control.tint[2] ),
    .B(\pll_control.tint[3] ),
    .C(\pll_control.tint[4] ),
    .ZN(_254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _509_ (.A1(net2),
    .A2(net20),
    .ZN(_255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _510_ (.A1(_254_),
    .A2(net2),
    .B(_255_),
    .ZN(\itrim[20] ));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _511_ (.A1(_223_),
    .A2(_126_),
    .A3(\pll_control.tint[0] ),
    .Z(_256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _512_ (.A1(net2),
    .A2(net21),
    .ZN(_257_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _513_ (.A1(_243_),
    .A2(_256_),
    .B(_257_),
    .ZN(\itrim[21] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _514_ (.A1(_234_),
    .A2(_214_),
    .ZN(_258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _515_ (.A1(net2),
    .A2(net22),
    .ZN(_259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _516_ (.A1(_258_),
    .A2(_259_),
    .ZN(\itrim[22] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _517_ (.I0(\pll_control.tint[4] ),
    .I1(net23),
    .S(net2),
    .Z(\itrim[23] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _518_ (.I0(_110_),
    .I1(net24),
    .S(net2),
    .Z(\itrim[24] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _519_ (.A1(net2),
    .A2(net25),
    .ZN(_260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _520_ (.A1(_240_),
    .A2(_209_),
    .B(_260_),
    .ZN(\itrim[25] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _521_ (.A1(_120_),
    .A2(_123_),
    .ZN(_261_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _522_ (.I0(_261_),
    .I1(net26),
    .S(net2),
    .Z(\itrim[2] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _523_ (.I0(_124_),
    .I1(net27),
    .S(net2),
    .Z(\itrim[3] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _524_ (.A1(net2),
    .A2(net28),
    .ZN(_262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _525_ (.A1(_203_),
    .A2(_262_),
    .ZN(\itrim[4] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _526_ (.A1(net2),
    .A2(net29),
    .ZN(_263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _527_ (.A1(_251_),
    .A2(_263_),
    .ZN(\itrim[5] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _528_ (.I(_124_),
    .ZN(_264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _529_ (.A1(_264_),
    .A2(_126_),
    .ZN(_265_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _530_ (.I0(_265_),
    .I1(net30),
    .S(net2),
    .Z(\itrim[6] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _531_ (.A1(net2),
    .A2(net31),
    .ZN(_266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _532_ (.A1(_219_),
    .A2(_266_),
    .ZN(\itrim[7] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _533_ (.A1(net2),
    .A2(net32),
    .ZN(_267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _534_ (.A1(_209_),
    .A2(_267_),
    .ZN(\itrim[8] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _535_ (.A1(net2),
    .A2(net33),
    .ZN(_268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _536_ (.A1(_213_),
    .A2(_268_),
    .ZN(\itrim[9] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input26 (.I(ext_trim[3]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count0[0]$_DFFE_PP0P_  (.D(_048_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.count0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count0[1]$_DFFE_PP0P_  (.D(_049_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.count0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count0[2]$_DFFE_PP0P_  (.D(_050_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.count0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count0[3]$_DFFE_PP0P_  (.D(_051_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.count0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count0[4]$_DFFE_PP0P_  (.D(_052_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.count0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count1[0]$_DFFE_PP0N_  (.D(_053_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.count1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count1[1]$_DFFE_PP0N_  (.D(_054_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.count1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count1[2]$_DFFE_PP0N_  (.D(_055_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.count1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count1[3]$_DFFE_PP0N_  (.D(_056_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.count1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count1[4]$_DFFE_PP0N_  (.D(_057_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.count1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.oscbuf[0]$_DFF_PP0_  (.D(osc),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.oscbuf[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.oscbuf[1]$_DFF_PP0_  (.D(\pll_control.oscbuf[0] ),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.oscbuf[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.oscbuf[2]$_DFF_PP0_  (.D(\pll_control.oscbuf[1] ),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.oscbuf[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.prep[0]$_DFFE_PP0N_  (.D(_058_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.prep[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.prep[1]$_DFFE_PP0N_  (.D(_059_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.prep[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.prep[2]$_DFFE_PP0N_  (.D(_060_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.prep[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.tval[0]$_DFFE_PP0P_  (.D(_061_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.tval[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.tval[1]$_DFFE_PP0P_  (.D(_062_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.tval[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.tval[2]$_DFFE_PP0P_  (.D(_063_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.tint[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.tval[3]$_DFFE_PP0P_  (.D(_064_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.tint[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.tval[4]$_DFFE_PP0P_  (.D(_065_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.tint[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.tval[5]$_DFFE_PP0P_  (.D(_066_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.tint[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.tval[6]$_DFFE_PP0P_  (.D(_067_),
    .RN(_047_),
    .CLK(net35),
    .Q(\pll_control.tint[4] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input25 (.I(ext_trim[2]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input24 (.I(ext_trim[25]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[0].id.delayen0  (.EN(\itrim[0] ),
    .I(\ringosc.dstage[0].id.d2 ),
    .ZN(\ringosc.dstage[0].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[0].id.delayen1  (.EN(\itrim[13] ),
    .I(\ringosc.dstage[0].id.in ),
    .ZN(\ringosc.dstage[0].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[0].id.delayenb0  (.EN(\ringosc.dstage[0].id.trim0b ),
    .I(\ringosc.dstage[0].id.in ),
    .ZN(\ringosc.dstage[0].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[0].id.delayenb1  (.EN(\ringosc.dstage[0].id.trim1b ),
    .I(\ringosc.dstage[0].id.in ),
    .ZN(\ringosc.dstage[0].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[0].id.delayint0  (.I(\ringosc.dstage[0].id.d1 ),
    .ZN(\ringosc.dstage[0].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[0].id.trim0bar  (.I(\itrim[0] ),
    .ZN(\ringosc.dstage[0].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[0].id.trim1bar  (.I(\itrim[13] ),
    .ZN(\ringosc.dstage[0].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input23 (.I(ext_trim[24]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input22 (.I(ext_trim[23]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[10].id.delayen0  (.EN(\itrim[10] ),
    .I(\ringosc.dstage[10].id.d2 ),
    .ZN(\ringosc.dstage[10].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[10].id.delayen1  (.EN(\itrim[23] ),
    .I(\ringosc.dstage[10].id.in ),
    .ZN(\ringosc.dstage[10].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[10].id.delayenb0  (.EN(\ringosc.dstage[10].id.trim0b ),
    .I(\ringosc.dstage[10].id.in ),
    .ZN(\ringosc.dstage[10].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[10].id.delayenb1  (.EN(\ringosc.dstage[10].id.trim1b ),
    .I(\ringosc.dstage[10].id.in ),
    .ZN(\ringosc.dstage[10].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[10].id.delayint0  (.I(\ringosc.dstage[10].id.d1 ),
    .ZN(\ringosc.dstage[10].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[10].id.trim0bar  (.I(\itrim[10] ),
    .ZN(\ringosc.dstage[10].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[10].id.trim1bar  (.I(\itrim[23] ),
    .ZN(\ringosc.dstage[10].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input21 (.I(ext_trim[22]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input20 (.I(ext_trim[21]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[11].id.delayen0  (.EN(\itrim[11] ),
    .I(\ringosc.dstage[11].id.d2 ),
    .ZN(\ringosc.dstage[11].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[11].id.delayen1  (.EN(\itrim[24] ),
    .I(\ringosc.dstage[10].id.out ),
    .ZN(\ringosc.dstage[11].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[11].id.delayenb0  (.EN(\ringosc.dstage[11].id.trim0b ),
    .I(\ringosc.dstage[10].id.out ),
    .ZN(\ringosc.dstage[11].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[11].id.delayenb1  (.EN(\ringosc.dstage[11].id.trim1b ),
    .I(\ringosc.dstage[10].id.out ),
    .ZN(\ringosc.dstage[11].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[11].id.delayint0  (.I(\ringosc.dstage[11].id.d1 ),
    .ZN(\ringosc.dstage[11].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[11].id.trim0bar  (.I(\itrim[11] ),
    .ZN(\ringosc.dstage[11].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[11].id.trim1bar  (.I(\itrim[24] ),
    .ZN(\ringosc.dstage[11].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input19 (.I(ext_trim[20]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input18 (.I(ext_trim[1]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[1].id.delayen0  (.EN(\itrim[1] ),
    .I(\ringosc.dstage[1].id.d2 ),
    .ZN(\ringosc.dstage[1].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[1].id.delayen1  (.EN(\itrim[14] ),
    .I(\ringosc.dstage[0].id.out ),
    .ZN(\ringosc.dstage[1].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[1].id.delayenb0  (.EN(\ringosc.dstage[1].id.trim0b ),
    .I(\ringosc.dstage[0].id.out ),
    .ZN(\ringosc.dstage[1].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[1].id.delayenb1  (.EN(\ringosc.dstage[1].id.trim1b ),
    .I(\ringosc.dstage[0].id.out ),
    .ZN(\ringosc.dstage[1].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[1].id.delayint0  (.I(\ringosc.dstage[1].id.d1 ),
    .ZN(\ringosc.dstage[1].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[1].id.trim0bar  (.I(\itrim[1] ),
    .ZN(\ringosc.dstage[1].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[1].id.trim1bar  (.I(\itrim[14] ),
    .ZN(\ringosc.dstage[1].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input17 (.I(ext_trim[19]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input16 (.I(ext_trim[18]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[2].id.delayen0  (.EN(\itrim[2] ),
    .I(\ringosc.dstage[2].id.d2 ),
    .ZN(\ringosc.dstage[2].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[2].id.delayen1  (.EN(\itrim[15] ),
    .I(\ringosc.dstage[1].id.out ),
    .ZN(\ringosc.dstage[2].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[2].id.delayenb0  (.EN(\ringosc.dstage[2].id.trim0b ),
    .I(\ringosc.dstage[1].id.out ),
    .ZN(\ringosc.dstage[2].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[2].id.delayenb1  (.EN(\ringosc.dstage[2].id.trim1b ),
    .I(\ringosc.dstage[1].id.out ),
    .ZN(\ringosc.dstage[2].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[2].id.delayint0  (.I(\ringosc.dstage[2].id.d1 ),
    .ZN(\ringosc.dstage[2].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[2].id.trim0bar  (.I(\itrim[2] ),
    .ZN(\ringosc.dstage[2].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[2].id.trim1bar  (.I(\itrim[15] ),
    .ZN(\ringosc.dstage[2].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input15 (.I(ext_trim[17]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input14 (.I(ext_trim[16]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[3].id.delayen0  (.EN(\itrim[3] ),
    .I(\ringosc.dstage[3].id.d2 ),
    .ZN(\ringosc.dstage[3].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[3].id.delayen1  (.EN(\itrim[16] ),
    .I(\ringosc.dstage[2].id.out ),
    .ZN(\ringosc.dstage[3].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[3].id.delayenb0  (.EN(\ringosc.dstage[3].id.trim0b ),
    .I(\ringosc.dstage[2].id.out ),
    .ZN(\ringosc.dstage[3].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[3].id.delayenb1  (.EN(\ringosc.dstage[3].id.trim1b ),
    .I(\ringosc.dstage[2].id.out ),
    .ZN(\ringosc.dstage[3].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[3].id.delayint0  (.I(\ringosc.dstage[3].id.d1 ),
    .ZN(\ringosc.dstage[3].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[3].id.trim0bar  (.I(\itrim[3] ),
    .ZN(\ringosc.dstage[3].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[3].id.trim1bar  (.I(\itrim[16] ),
    .ZN(\ringosc.dstage[3].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input13 (.I(ext_trim[15]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input12 (.I(ext_trim[14]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[4].id.delayen0  (.EN(\itrim[4] ),
    .I(\ringosc.dstage[4].id.d2 ),
    .ZN(\ringosc.dstage[4].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[4].id.delayen1  (.EN(\itrim[17] ),
    .I(\ringosc.dstage[3].id.out ),
    .ZN(\ringosc.dstage[4].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[4].id.delayenb0  (.EN(\ringosc.dstage[4].id.trim0b ),
    .I(\ringosc.dstage[3].id.out ),
    .ZN(\ringosc.dstage[4].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[4].id.delayenb1  (.EN(\ringosc.dstage[4].id.trim1b ),
    .I(\ringosc.dstage[3].id.out ),
    .ZN(\ringosc.dstage[4].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[4].id.delayint0  (.I(\ringosc.dstage[4].id.d1 ),
    .ZN(\ringosc.dstage[4].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[4].id.trim0bar  (.I(\itrim[4] ),
    .ZN(\ringosc.dstage[4].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[4].id.trim1bar  (.I(\itrim[17] ),
    .ZN(\ringosc.dstage[4].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input11 (.I(ext_trim[13]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input10 (.I(ext_trim[12]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[5].id.delayen0  (.EN(\itrim[5] ),
    .I(\ringosc.dstage[5].id.d2 ),
    .ZN(\ringosc.dstage[5].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[5].id.delayen1  (.EN(\itrim[18] ),
    .I(\ringosc.dstage[4].id.out ),
    .ZN(\ringosc.dstage[5].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[5].id.delayenb0  (.EN(\ringosc.dstage[5].id.trim0b ),
    .I(\ringosc.dstage[4].id.out ),
    .ZN(\ringosc.dstage[5].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[5].id.delayenb1  (.EN(\ringosc.dstage[5].id.trim1b ),
    .I(\ringosc.dstage[4].id.out ),
    .ZN(\ringosc.dstage[5].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[5].id.delayint0  (.I(\ringosc.dstage[5].id.d1 ),
    .ZN(\ringosc.dstage[5].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[5].id.trim0bar  (.I(\itrim[5] ),
    .ZN(\ringosc.dstage[5].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[5].id.trim1bar  (.I(\itrim[18] ),
    .ZN(\ringosc.dstage[5].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input9 (.I(ext_trim[11]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input8 (.I(ext_trim[10]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[6].id.delayen0  (.EN(\itrim[6] ),
    .I(\ringosc.dstage[6].id.d2 ),
    .ZN(\ringosc.dstage[6].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[6].id.delayen1  (.EN(\itrim[19] ),
    .I(\ringosc.dstage[5].id.out ),
    .ZN(\ringosc.dstage[6].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[6].id.delayenb0  (.EN(\ringosc.dstage[6].id.trim0b ),
    .I(\ringosc.dstage[5].id.out ),
    .ZN(\ringosc.dstage[6].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[6].id.delayenb1  (.EN(\ringosc.dstage[6].id.trim1b ),
    .I(\ringosc.dstage[5].id.out ),
    .ZN(\ringosc.dstage[6].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[6].id.delayint0  (.I(\ringosc.dstage[6].id.d1 ),
    .ZN(\ringosc.dstage[6].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[6].id.trim0bar  (.I(\itrim[6] ),
    .ZN(\ringosc.dstage[6].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[6].id.trim1bar  (.I(\itrim[19] ),
    .ZN(\ringosc.dstage[6].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input7 (.I(ext_trim[0]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input6 (.I(enable),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[7].id.delayen0  (.EN(\itrim[7] ),
    .I(\ringosc.dstage[7].id.d2 ),
    .ZN(\ringosc.dstage[7].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[7].id.delayen1  (.EN(\itrim[20] ),
    .I(\ringosc.dstage[6].id.out ),
    .ZN(\ringosc.dstage[7].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[7].id.delayenb0  (.EN(\ringosc.dstage[7].id.trim0b ),
    .I(\ringosc.dstage[6].id.out ),
    .ZN(\ringosc.dstage[7].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[7].id.delayenb1  (.EN(\ringosc.dstage[7].id.trim1b ),
    .I(\ringosc.dstage[6].id.out ),
    .ZN(\ringosc.dstage[7].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[7].id.delayint0  (.I(\ringosc.dstage[7].id.d1 ),
    .ZN(\ringosc.dstage[7].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[7].id.trim0bar  (.I(\itrim[7] ),
    .ZN(\ringosc.dstage[7].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[7].id.trim1bar  (.I(\itrim[20] ),
    .ZN(\ringosc.dstage[7].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input5 (.I(div[4]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input4 (.I(div[3]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[8].id.delayen0  (.EN(\itrim[8] ),
    .I(\ringosc.dstage[8].id.d2 ),
    .ZN(\ringosc.dstage[8].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[8].id.delayen1  (.EN(\itrim[21] ),
    .I(\ringosc.dstage[7].id.out ),
    .ZN(\ringosc.dstage[8].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[8].id.delayenb0  (.EN(\ringosc.dstage[8].id.trim0b ),
    .I(\ringosc.dstage[7].id.out ),
    .ZN(\ringosc.dstage[8].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[8].id.delayenb1  (.EN(\ringosc.dstage[8].id.trim1b ),
    .I(\ringosc.dstage[7].id.out ),
    .ZN(\ringosc.dstage[8].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[8].id.delayint0  (.I(\ringosc.dstage[8].id.d1 ),
    .ZN(\ringosc.dstage[8].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[8].id.trim0bar  (.I(\itrim[8] ),
    .ZN(\ringosc.dstage[8].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[8].id.trim1bar  (.I(\itrim[21] ),
    .ZN(\ringosc.dstage[8].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input3 (.I(div[2]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input2 (.I(div[1]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[9].id.delayen0  (.EN(\itrim[9] ),
    .I(\ringosc.dstage[9].id.d2 ),
    .ZN(\ringosc.dstage[10].id.in ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[9].id.delayen1  (.EN(\itrim[22] ),
    .I(\ringosc.dstage[8].id.out ),
    .ZN(\ringosc.dstage[9].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[9].id.delayenb0  (.EN(\ringosc.dstage[9].id.trim0b ),
    .I(\ringosc.dstage[8].id.out ),
    .ZN(\ringosc.dstage[10].id.in ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[9].id.delayenb1  (.EN(\ringosc.dstage[9].id.trim1b ),
    .I(\ringosc.dstage[8].id.out ),
    .ZN(\ringosc.dstage[9].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[9].id.delayint0  (.I(\ringosc.dstage[9].id.d1 ),
    .ZN(\ringosc.dstage[9].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[9].id.trim0bar  (.I(\itrim[9] ),
    .ZN(\ringosc.dstage[9].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[9].id.trim1bar  (.I(\itrim[22] ),
    .ZN(\ringosc.dstage[9].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 \ringosc.ibufp00  (.I(\ringosc.dstage[0].id.in ),
    .ZN(\ringosc.c[0] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_8 \ringosc.ibufp01  (.I(\ringosc.c[0] ),
    .ZN(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.ibufp10  (.I(\ringosc.dstage[5].id.out ),
    .ZN(\ringosc.c[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.ibufp11  (.I(\ringosc.c[1] ),
    .ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 \ringosc.iss.ctrlen0  (.A1(ireset),
    .A2(\itrim[12] ),
    .ZN(\ringosc.iss.ctrl0b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 input1 (.I(dco),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.iss.delayen0  (.EN(\itrim[12] ),
    .I(\ringosc.iss.d2 ),
    .ZN(\ringosc.dstage[0].id.in ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.iss.delayen1  (.EN(\itrim[25] ),
    .I(\ringosc.dstage[11].id.out ),
    .ZN(\ringosc.iss.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.iss.delayenb0  (.EN(\ringosc.iss.ctrl0b ),
    .I(\ringosc.dstage[11].id.out ),
    .ZN(\ringosc.dstage[0].id.in ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.iss.delayenb1  (.EN(\ringosc.iss.trim1b ),
    .I(\ringosc.dstage[11].id.out ),
    .ZN(\ringosc.iss.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.iss.delayint0  (.I(\ringosc.iss.d1 ),
    .ZN(\ringosc.iss.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.iss.reseten0  (.EN(ireset),
    .I(net1),
    .ZN(\ringosc.dstage[0].id.in ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.iss.trim1bar  (.I(\itrim[25] ),
    .ZN(\ringosc.iss.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__tieh \ringosc.iss.reseten0_1  (.Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_184 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input33 (.I(resetb),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output34 (.I(net35),
    .Z(clockp[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output35 (.I(net36),
    .Z(clockp[1]));
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_0_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_0_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_0_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_0_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_1_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_1_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_1_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_1_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_1_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_2_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_2_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_2_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_2_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_2_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_2_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_2_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_2_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_2_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_2_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_2_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_2_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_2_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_3_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_3_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_3_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_3_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_3_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_3_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_3_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_3_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_3_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_3_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_3_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_3_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_3_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_3_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_4_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_4_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_4_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_4_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_4_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_4_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_4_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_4_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_4_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_4_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_4_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_6_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_6_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_6_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_6_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_6_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_6_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_7_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_7_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_7_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_7_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_7_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_7_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_8_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_8_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_8_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_8_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_8_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_9_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_9_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_9_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_9_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_10_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_10_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_10_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_10_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_10_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_10_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_10_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_10_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_10_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_10_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_11_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_11_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_11_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_11_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_11_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_11_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_11_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_11_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_12_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_12_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_12_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_12_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_12_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_13_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_13_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_14_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_14_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_14_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_14_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_14_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_15_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_15_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_16_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_16_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_16_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_16_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_16_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_16_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_16_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_16_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_16_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_16_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_16_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_17_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_17_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_17_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_17_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_17_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_17_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_17_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_17_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_18_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_18_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_18_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_18_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_18_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_18_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_18_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_18_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_18_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_18_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_19_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_19_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_19_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_19_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_19_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_19_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_19_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_20_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_20_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_20_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_20_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_20_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_20_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_20_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_20_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_20_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_20_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_21_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_21_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_21_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_21_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_21_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_21_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_21_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_21_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_22_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_22_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_22_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_22_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_22_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_22_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_22_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_22_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_22_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_22_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_22_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_22_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_23_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_23_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_23_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_23_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_23_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_23_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_23_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_23_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_23_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_23_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_23_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_23_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_23_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_24_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_24_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_24_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_24_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_24_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_24_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_25_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_25_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_25_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_25_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_25_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_25_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_25_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_25_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_25_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_25_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_25_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_25_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_25_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_25_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_25_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_26_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_26_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_26_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_26_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_26_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_26_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_26_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_26_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_26_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_27_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_27_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_27_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_27_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_27_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_27_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_27_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_27_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_27_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_27_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_27_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_27_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_28_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_28_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_28_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_28_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_28_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_28_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_28_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_28_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_28_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_28_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_28_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_28_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_29_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_29_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_29_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_29_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_29_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_29_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_29_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_29_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_29_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_29_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_29_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_30_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_30_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_30_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_30_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_30_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_30_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_30_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_30_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_30_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_31_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_31_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_31_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_31_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_31_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_31_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_31_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_31_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_31_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_31_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_31_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_31_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_32_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_32_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_32_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_32_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_32_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_32_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_32_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_32_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_32_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_32_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_32_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_32_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_32_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_33_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_33_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_33_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_33_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_33_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_33_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_33_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_33_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_33_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_33_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_33_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_33_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_33_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_33_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_34_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_34_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_34_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_34_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_34_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_34_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_34_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_34_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_35_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_35_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_35_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_35_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_35_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_36_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_36_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_36_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_36_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_36_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_36_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_36_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_36_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_37_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_37_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_37_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_37_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_37_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_37_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_37_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_37_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_37_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_37_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_37_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_37_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_38_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_38_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_38_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_38_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_38_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_38_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_39_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_39_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_39_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_39_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_39_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_39_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_39_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_39_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_40_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_40_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_40_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_40_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_40_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_40_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_40_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_40_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_40_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_41_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_41_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_41_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_41_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_41_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_41_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_41_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_41_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_41_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_42_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_42_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_42_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_42_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_42_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_42_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_43_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_43_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_43_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_43_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_43_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_43_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_43_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_43_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_43_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_44_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_44_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_44_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_44_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_44_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_44_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_44_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_44_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_45_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_45_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_45_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_45_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_45_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_45_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_45_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_45_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_45_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_45_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_45_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_45_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_46_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_46_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_46_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_46_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_46_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_46_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_46_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_46_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_46_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_47_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_47_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_47_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_47_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_47_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_47_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_47_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_47_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_47_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_48_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_48_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_48_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_48_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_48_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_48_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_48_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_48_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_48_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_48_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_49_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_49_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_49_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_49_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_49_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_49_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_49_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_50_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_50_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_50_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_50_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_50_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_50_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_50_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_50_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_51_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_51_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_51_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_51_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_51_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_51_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_51_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_51_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_51_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_52_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_52_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_52_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_52_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_52_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_52_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_52_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_52_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_52_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_52_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_52_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_53_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_53_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_53_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_53_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_53_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_53_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_53_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_54_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_54_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_54_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_54_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_54_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_54_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_54_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_54_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_55_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_55_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_55_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_55_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_55_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_55_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_55_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_55_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_55_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_56_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_56_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_56_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_56_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_56_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_56_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_56_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_57_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_57_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_57_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_57_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_57_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_57_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_57_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_57_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_57_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_57_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_57_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_57_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_57_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_58_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_58_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_58_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_58_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_58_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_58_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_58_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_58_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_58_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_58_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_58_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_58_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_59_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_59_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_59_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_59_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_59_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_59_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_59_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_59_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_59_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_59_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_60_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_60_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_60_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_60_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_60_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_60_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_60_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_60_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_60_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_60_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_60_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_60_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_432 ();
endmodule
