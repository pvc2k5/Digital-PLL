module digital_pll (dco,
    enable,
    osc,
    resetb,
    clockp,
    div,
    ext_trim);
 input dco;
 input enable;
 input osc;
 input resetb;
 output [1:0] clockp;
 input [4:0] div;
 input [25:0] ext_trim;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire net33;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire net32;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire net31;
 wire _167_;
 wire net30;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire net29;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire net28;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire net36;
 wire net37;
 wire ireset;
 wire \itrim[0] ;
 wire \itrim[10] ;
 wire \itrim[11] ;
 wire \itrim[12] ;
 wire \itrim[13] ;
 wire \itrim[14] ;
 wire \itrim[15] ;
 wire \itrim[16] ;
 wire \itrim[17] ;
 wire \itrim[18] ;
 wire \itrim[19] ;
 wire \itrim[1] ;
 wire \itrim[20] ;
 wire \itrim[21] ;
 wire \itrim[22] ;
 wire \itrim[23] ;
 wire \itrim[24] ;
 wire \itrim[25] ;
 wire \itrim[2] ;
 wire \itrim[3] ;
 wire \itrim[4] ;
 wire \itrim[5] ;
 wire \itrim[6] ;
 wire \itrim[7] ;
 wire \itrim[8] ;
 wire \itrim[9] ;
 wire net27;
 wire \pll_control.count0[0] ;
 wire \pll_control.count0[1] ;
 wire \pll_control.count0[2] ;
 wire \pll_control.count0[3] ;
 wire \pll_control.count0[4] ;
 wire \pll_control.count1[0] ;
 wire \pll_control.count1[1] ;
 wire \pll_control.count1[2] ;
 wire \pll_control.count1[3] ;
 wire \pll_control.count1[4] ;
 wire \pll_control.oscbuf[0] ;
 wire \pll_control.oscbuf[1] ;
 wire \pll_control.oscbuf[2] ;
 wire \pll_control.prep[0] ;
 wire \pll_control.prep[1] ;
 wire \pll_control.prep[2] ;
 wire \pll_control.tint[0] ;
 wire \pll_control.tint[1] ;
 wire \pll_control.tint[2] ;
 wire \pll_control.tint[3] ;
 wire \pll_control.tint[4] ;
 wire \pll_control.tval[0] ;
 wire \pll_control.tval[1] ;
 wire \ringosc.c[0] ;
 wire \ringosc.c[1] ;
 wire net25;
 wire \ringosc.dstage[0].id.d1 ;
 wire \ringosc.dstage[0].id.d2 ;
 wire \ringosc.dstage[0].id.in ;
 wire \ringosc.dstage[0].id.out ;
 wire \ringosc.dstage[0].id.trim0b ;
 wire \ringosc.dstage[0].id.trim1b ;
 wire net26;
 wire net23;
 wire \ringosc.dstage[10].id.d1 ;
 wire \ringosc.dstage[10].id.d2 ;
 wire \ringosc.dstage[10].id.in ;
 wire \ringosc.dstage[10].id.out ;
 wire \ringosc.dstage[10].id.trim0b ;
 wire \ringosc.dstage[10].id.trim1b ;
 wire net24;
 wire net21;
 wire \ringosc.dstage[11].id.d1 ;
 wire \ringosc.dstage[11].id.d2 ;
 wire \ringosc.dstage[11].id.out ;
 wire \ringosc.dstage[11].id.trim0b ;
 wire \ringosc.dstage[11].id.trim1b ;
 wire net22;
 wire net19;
 wire \ringosc.dstage[1].id.d1 ;
 wire \ringosc.dstage[1].id.d2 ;
 wire \ringosc.dstage[1].id.out ;
 wire \ringosc.dstage[1].id.trim0b ;
 wire \ringosc.dstage[1].id.trim1b ;
 wire net20;
 wire net17;
 wire \ringosc.dstage[2].id.d1 ;
 wire \ringosc.dstage[2].id.d2 ;
 wire \ringosc.dstage[2].id.out ;
 wire \ringosc.dstage[2].id.trim0b ;
 wire \ringosc.dstage[2].id.trim1b ;
 wire net18;
 wire net15;
 wire \ringosc.dstage[3].id.d1 ;
 wire \ringosc.dstage[3].id.d2 ;
 wire \ringosc.dstage[3].id.out ;
 wire \ringosc.dstage[3].id.trim0b ;
 wire \ringosc.dstage[3].id.trim1b ;
 wire net16;
 wire net13;
 wire \ringosc.dstage[4].id.d1 ;
 wire \ringosc.dstage[4].id.d2 ;
 wire \ringosc.dstage[4].id.out ;
 wire \ringosc.dstage[4].id.trim0b ;
 wire \ringosc.dstage[4].id.trim1b ;
 wire net14;
 wire net11;
 wire \ringosc.dstage[5].id.d1 ;
 wire \ringosc.dstage[5].id.d2 ;
 wire \ringosc.dstage[5].id.out ;
 wire \ringosc.dstage[5].id.trim0b ;
 wire \ringosc.dstage[5].id.trim1b ;
 wire net12;
 wire net9;
 wire \ringosc.dstage[6].id.d1 ;
 wire \ringosc.dstage[6].id.d2 ;
 wire \ringosc.dstage[6].id.out ;
 wire \ringosc.dstage[6].id.trim0b ;
 wire \ringosc.dstage[6].id.trim1b ;
 wire net10;
 wire net7;
 wire \ringosc.dstage[7].id.d1 ;
 wire \ringosc.dstage[7].id.d2 ;
 wire \ringosc.dstage[7].id.out ;
 wire \ringosc.dstage[7].id.trim0b ;
 wire \ringosc.dstage[7].id.trim1b ;
 wire net8;
 wire net5;
 wire \ringosc.dstage[8].id.d1 ;
 wire \ringosc.dstage[8].id.d2 ;
 wire \ringosc.dstage[8].id.out ;
 wire \ringosc.dstage[8].id.trim0b ;
 wire \ringosc.dstage[8].id.trim1b ;
 wire net6;
 wire net3;
 wire \ringosc.dstage[9].id.d1 ;
 wire \ringosc.dstage[9].id.d2 ;
 wire \ringosc.dstage[9].id.trim0b ;
 wire \ringosc.dstage[9].id.trim1b ;
 wire net4;
 wire \ringosc.iss.ctrl0b ;
 wire net2;
 wire \ringosc.iss.d1 ;
 wire \ringosc.iss.d2 ;
 wire \ringosc.iss.trim1b ;
 wire net1;
 wire net34;
 wire net35;

 gf180mcu_fd_sc_mcu7t5v0__and3_2 _274_ (.A1(\pll_control.count0[2] ),
    .A2(\pll_control.count0[3] ),
    .A3(_032_),
    .Z(_034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _275_ (.A1(net8),
    .A2(net35),
    .ZN(ireset));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input32 (.I(ext_trim[8]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _277_ (.A1(ireset),
    .A2(net2),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _278_ (.I(net7),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _279_ (.I(_006_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _280_ (.A1(_001_),
    .A2(_010_),
    .B(_009_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _281_ (.I(_008_),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _282_ (.I(_007_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _283_ (.A1(_070_),
    .A2(_071_),
    .B(_072_),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _284_ (.A1(_069_),
    .A2(_073_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _285_ (.I(net6),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _286_ (.I(net5),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _287_ (.I(net4),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _288_ (.A1(_023_),
    .A2(_020_),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _289_ (.I(_019_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _290_ (.A1(_074_),
    .A2(_075_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _291_ (.A1(_076_),
    .A2(_016_),
    .B(_015_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _292_ (.I(_030_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _293_ (.A1(_078_),
    .A2(_027_),
    .B(_026_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _294_ (.A1(_016_),
    .A2(_020_),
    .A3(_024_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _295_ (.A1(_079_),
    .A2(_080_),
    .Z(_081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _296_ (.A1(_077_),
    .A2(_081_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _297_ (.A1(_027_),
    .A2(_031_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _298_ (.A1(_080_),
    .A2(_083_),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _299_ (.I(_084_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _300_ (.A1(_082_),
    .A2(_085_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _301_ (.A1(_010_),
    .A2(_011_),
    .B(_009_),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _302_ (.A1(_000_),
    .A2(_010_),
    .A3(_012_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _303_ (.A1(_087_),
    .A2(_088_),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _304_ (.A1(_006_),
    .A2(_008_),
    .Z(_090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _305_ (.A1(_089_),
    .A2(_090_),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _306_ (.A1(_006_),
    .A2(_007_),
    .Z(_092_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _307_ (.A1(_092_),
    .A2(_005_),
    .Z(_093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _308_ (.I(_093_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _309_ (.A1(_091_),
    .A2(_094_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _310_ (.I(_095_),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _311_ (.A1(_086_),
    .A2(_096_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _312_ (.A1(_071_),
    .A2(_089_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _313_ (.A1(_001_),
    .A2(_010_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _314_ (.I(_028_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _315_ (.I(_035_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _316_ (.A1(\pll_control.count0[0] ),
    .A2(_097_),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _317_ (.I(\pll_control.oscbuf[1] ),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _318_ (.A1(_099_),
    .A2(\pll_control.oscbuf[2] ),
    .Z(_100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _319_ (.A1(_099_),
    .A2(\pll_control.oscbuf[2] ),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _320_ (.A1(_100_),
    .A2(_101_),
    .Z(_102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input31 (.I(ext_trim[7]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _322_ (.A1(_098_),
    .A2(_102_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _323_ (.I0(_033_),
    .I1(\pll_control.count0[1] ),
    .S(_035_),
    .Z(_104_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _324_ (.A1(_104_),
    .A2(_102_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _325_ (.I(_102_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _326_ (.A1(_097_),
    .A2(_032_),
    .B(\pll_control.count0[2] ),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _327_ (.A1(_097_),
    .A2(\pll_control.count0[2] ),
    .A3(_032_),
    .Z(_107_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _328_ (.A1(_105_),
    .A2(_106_),
    .A3(_107_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _329_ (.A1(_097_),
    .A2(\pll_control.count0[2] ),
    .A3(\pll_control.count0[0] ),
    .A4(\pll_control.count0[1] ),
    .Z(_108_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _330_ (.A1(_108_),
    .A2(\pll_control.count0[3] ),
    .Z(_109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _331_ (.A1(_108_),
    .A2(\pll_control.count0[3] ),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _332_ (.A1(_109_),
    .A2(_102_),
    .A3(_110_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _333_ (.I0(_036_),
    .I1(\pll_control.count0[4] ),
    .S(_035_),
    .Z(_111_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _334_ (.A1(_111_),
    .A2(_102_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _335_ (.I(\pll_control.tint[3] ),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _336_ (.I(\pll_control.tint[2] ),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _337_ (.A1(_112_),
    .A2(_113_),
    .Z(_114_));
 gf180mcu_fd_sc_mcu7t5v0__inv_8 _338_ (.I(\pll_control.tint[4] ),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _339_ (.A1(_114_),
    .A2(_115_),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _340_ (.A1(\pll_control.tval[0] ),
    .A2(\pll_control.tval[1] ),
    .Z(_117_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _341_ (.I(\pll_control.tint[1] ),
    .ZN(_118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _342_ (.I(\pll_control.tint[0] ),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _343_ (.A1(_118_),
    .A2(_119_),
    .Z(_120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _344_ (.I(_120_),
    .ZN(_121_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _345_ (.A1(_116_),
    .A2(_117_),
    .A3(_121_),
    .Z(_122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _346_ (.I(_082_),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _347_ (.A1(_096_),
    .A2(_122_),
    .A3(_123_),
    .ZN(_124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _348_ (.A1(_124_),
    .A2(_002_),
    .ZN(_125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _349_ (.A1(_077_),
    .A2(_081_),
    .B(_084_),
    .ZN(_126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _350_ (.A1(\pll_control.tint[1] ),
    .A2(\pll_control.tint[0] ),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _351_ (.I(_127_),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _352_ (.A1(\pll_control.tint[3] ),
    .A2(\pll_control.tint[4] ),
    .Z(_129_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _353_ (.A1(\pll_control.tval[0] ),
    .A2(\pll_control.tval[1] ),
    .Z(_130_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _354_ (.A1(_128_),
    .A2(_129_),
    .A3(_130_),
    .A4(\pll_control.tint[2] ),
    .Z(_131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _355_ (.A1(_126_),
    .A2(_095_),
    .B(_131_),
    .ZN(_132_));
 gf180mcu_fd_sc_mcu7t5v0__and4_4 _356_ (.A1(_105_),
    .A2(\pll_control.prep[1] ),
    .A3(\pll_control.prep[0] ),
    .A4(\pll_control.prep[2] ),
    .Z(_133_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _357_ (.A1(_125_),
    .A2(_132_),
    .A3(_133_),
    .ZN(_134_));
 gf180mcu_fd_sc_mcu7t5v0__inv_8 _358_ (.I(_134_),
    .ZN(_135_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _359_ (.I(\pll_control.tval[0] ),
    .ZN(_136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _360_ (.A1(_135_),
    .A2(_136_),
    .ZN(_137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _361_ (.A1(_134_),
    .A2(\pll_control.tval[0] ),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _362_ (.A1(_137_),
    .A2(_138_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _363_ (.A1(_135_),
    .A2(_004_),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _364_ (.A1(_134_),
    .A2(\pll_control.tval[1] ),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _365_ (.A1(_139_),
    .A2(_140_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _366_ (.I(_040_),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _367_ (.A1(_003_),
    .A2(_141_),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _368_ (.A1(_135_),
    .A2(_142_),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _369_ (.A1(_134_),
    .A2(\pll_control.tint[0] ),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _370_ (.A1(_143_),
    .A2(_144_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _371_ (.I(_042_),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _372_ (.I(_038_),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _373_ (.A1(_040_),
    .A2(_037_),
    .B(_039_),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _374_ (.A1(_136_),
    .A2(_146_),
    .A3(_141_),
    .B(_147_),
    .ZN(_148_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _375_ (.A1(_145_),
    .A2(_148_),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _376_ (.A1(_135_),
    .A2(_149_),
    .ZN(_150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _377_ (.A1(_134_),
    .A2(\pll_control.tint[1] ),
    .ZN(_151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _378_ (.A1(_150_),
    .A2(_151_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _379_ (.I(_044_),
    .ZN(_152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _380_ (.I(_003_),
    .ZN(_153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _381_ (.A1(_042_),
    .A2(_039_),
    .B(_041_),
    .ZN(_154_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _382_ (.A1(_153_),
    .A2(_141_),
    .A3(_145_),
    .B(_154_),
    .ZN(_155_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _383_ (.A1(_152_),
    .A2(_155_),
    .ZN(_156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _384_ (.A1(_135_),
    .A2(_156_),
    .ZN(_157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _385_ (.A1(_134_),
    .A2(\pll_control.tint[2] ),
    .ZN(_158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _386_ (.A1(_157_),
    .A2(_158_),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _387_ (.A1(_042_),
    .A2(_044_),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _388_ (.A1(_159_),
    .A2(_146_),
    .A3(_141_),
    .Z(_160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _389_ (.A1(_044_),
    .A2(_041_),
    .B(_043_),
    .ZN(_161_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _390_ (.A1(_136_),
    .A2(_160_),
    .B1(_147_),
    .B2(_159_),
    .C(_161_),
    .ZN(_162_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _391_ (.A1(_046_),
    .A2(_162_),
    .Z(_163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _392_ (.A1(_135_),
    .A2(_163_),
    .ZN(_164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _393_ (.A1(_134_),
    .A2(\pll_control.tint[3] ),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _394_ (.A1(_164_),
    .A2(_165_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input30 (.I(ext_trim[6]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _396_ (.A1(_126_),
    .A2(_095_),
    .B(_115_),
    .ZN(_167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input29 (.I(ext_trim[5]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _398_ (.A1(_086_),
    .A2(\pll_control.tint[4] ),
    .A3(_096_),
    .ZN(_169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _399_ (.A1(_167_),
    .A2(_169_),
    .ZN(_170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _400_ (.A1(_044_),
    .A2(_046_),
    .ZN(_171_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _401_ (.A1(_171_),
    .A2(_153_),
    .A3(_141_),
    .A4(_145_),
    .Z(_172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _402_ (.A1(_046_),
    .A2(_043_),
    .B(_045_),
    .ZN(_173_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _403_ (.A1(_154_),
    .A2(_171_),
    .Z(_174_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _404_ (.A1(_172_),
    .A2(_173_),
    .A3(_174_),
    .Z(_175_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _405_ (.I(_175_),
    .ZN(_176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _406_ (.A1(_170_),
    .A2(_176_),
    .ZN(_177_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _407_ (.A1(_167_),
    .A2(_169_),
    .A3(_175_),
    .ZN(_178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _408_ (.A1(_177_),
    .A2(_178_),
    .ZN(_179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _409_ (.A1(_179_),
    .A2(_135_),
    .ZN(_180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _410_ (.A1(_134_),
    .A2(\pll_control.tint[4] ),
    .ZN(_181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _411_ (.A1(_180_),
    .A2(_181_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _412_ (.I0(\pll_control.count0[0] ),
    .I1(\pll_control.count1[0] ),
    .S(_102_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _413_ (.I0(\pll_control.count0[1] ),
    .I1(\pll_control.count1[1] ),
    .S(_102_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _414_ (.I0(\pll_control.count0[2] ),
    .I1(\pll_control.count1[2] ),
    .S(_102_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _415_ (.I0(\pll_control.count0[3] ),
    .I1(\pll_control.count1[3] ),
    .S(_102_),
    .Z(_056_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _416_ (.I0(\pll_control.count0[4] ),
    .I1(\pll_control.count1[4] ),
    .S(_102_),
    .Z(_057_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _417_ (.A1(_105_),
    .A2(\pll_control.prep[0] ),
    .Z(_058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _418_ (.I0(\pll_control.prep[0] ),
    .I1(\pll_control.prep[1] ),
    .S(_102_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _419_ (.I0(\pll_control.prep[1] ),
    .I1(\pll_control.prep[2] ),
    .S(_102_),
    .Z(_060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _420_ (.I(_116_),
    .ZN(_182_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _421_ (.A1(_182_),
    .A2(_120_),
    .Z(_183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input28 (.I(ext_trim[4]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _423_ (.A1(net2),
    .A2(net9),
    .ZN(_185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _424_ (.A1(_183_),
    .A2(net2),
    .B(_185_),
    .ZN(\itrim[0] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _425_ (.I(net2),
    .ZN(_186_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _426_ (.A1(_116_),
    .A2(_186_),
    .Z(_187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _427_ (.A1(_186_),
    .A2(_128_),
    .B(_187_),
    .ZN(_188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _428_ (.A1(net2),
    .A2(net10),
    .ZN(_189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _429_ (.A1(_188_),
    .A2(_189_),
    .ZN(\itrim[10] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _430_ (.A1(_112_),
    .A2(\pll_control.tint[2] ),
    .Z(_190_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _431_ (.A1(_190_),
    .A2(_128_),
    .Z(_191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _432_ (.A1(_191_),
    .A2(_115_),
    .ZN(_192_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _433_ (.A1(_120_),
    .A2(_190_),
    .Z(_193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _434_ (.A1(_193_),
    .A2(_115_),
    .ZN(_194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _435_ (.A1(_187_),
    .A2(_194_),
    .ZN(_195_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _436_ (.I(_195_),
    .ZN(_196_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _437_ (.A1(_115_),
    .A2(_119_),
    .A3(\pll_control.tint[1] ),
    .Z(_197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _438_ (.A1(_118_),
    .A2(\pll_control.tint[0] ),
    .ZN(_198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _439_ (.A1(_198_),
    .A2(\pll_control.tint[4] ),
    .ZN(_199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _440_ (.A1(_197_),
    .A2(_199_),
    .B(_190_),
    .ZN(_200_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _441_ (.A1(_196_),
    .A2(_200_),
    .Z(_201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _442_ (.A1(_113_),
    .A2(\pll_control.tint[3] ),
    .ZN(_202_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _443_ (.A1(_198_),
    .A2(_202_),
    .A3(\pll_control.tint[4] ),
    .Z(_203_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _444_ (.I(_202_),
    .ZN(_204_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _445_ (.A1(_120_),
    .A2(_204_),
    .A3(_115_),
    .Z(_205_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _446_ (.I(_205_),
    .ZN(_206_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _447_ (.A1(_192_),
    .A2(_201_),
    .A3(_203_),
    .A4(_206_),
    .ZN(_207_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _448_ (.A1(_197_),
    .A2(_204_),
    .Z(_208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _449_ (.A1(net2),
    .A2(net11),
    .ZN(_209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _450_ (.A1(_207_),
    .A2(_208_),
    .B(_209_),
    .ZN(\itrim[11] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _451_ (.A1(_199_),
    .A2(_190_),
    .Z(_210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _452_ (.A1(net2),
    .A2(net12),
    .ZN(_211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _453_ (.A1(_195_),
    .A2(_210_),
    .B(_211_),
    .ZN(\itrim[12] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _454_ (.A1(_206_),
    .A2(_192_),
    .Z(_212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _455_ (.A1(_201_),
    .A2(_212_),
    .ZN(_213_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _456_ (.A1(\pll_control.tint[3] ),
    .A2(\pll_control.tint[2] ),
    .Z(_214_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _457_ (.A1(_120_),
    .A2(_115_),
    .A3(_214_),
    .Z(_215_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _458_ (.A1(_204_),
    .A2(_115_),
    .A3(_128_),
    .Z(_216_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _459_ (.A1(_215_),
    .A2(_216_),
    .ZN(_217_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _460_ (.I(_208_),
    .ZN(_218_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _461_ (.A1(_217_),
    .A2(_218_),
    .A3(_203_),
    .ZN(_219_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _462_ (.A1(_213_),
    .A2(_219_),
    .Z(_220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _463_ (.A1(_199_),
    .A2(_214_),
    .ZN(_221_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _464_ (.I(_221_),
    .ZN(_222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _465_ (.A1(net2),
    .A2(net13),
    .ZN(_223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _466_ (.A1(_220_),
    .A2(_222_),
    .B(_223_),
    .ZN(\itrim[13] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _467_ (.A1(_114_),
    .A2(\pll_control.tint[4] ),
    .Z(_224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _468_ (.A1(_224_),
    .A2(_127_),
    .ZN(_225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _469_ (.A1(_128_),
    .A2(_214_),
    .ZN(_226_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _470_ (.A1(_226_),
    .A2(\pll_control.tint[4] ),
    .Z(_227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _471_ (.A1(_197_),
    .A2(_214_),
    .ZN(_228_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _472_ (.A1(_221_),
    .A2(_225_),
    .A3(_227_),
    .A4(_228_),
    .ZN(_229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _473_ (.A1(_229_),
    .A2(_219_),
    .ZN(_230_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _474_ (.A1(_114_),
    .A2(_128_),
    .Z(_231_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _475_ (.A1(_231_),
    .A2(\pll_control.tint[4] ),
    .Z(_232_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _476_ (.A1(_190_),
    .A2(\pll_control.tint[4] ),
    .A3(_118_),
    .Z(_233_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _477_ (.A1(_232_),
    .A2(_233_),
    .Z(_234_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _478_ (.I(_234_),
    .ZN(_235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _479_ (.A1(_230_),
    .A2(_235_),
    .ZN(_236_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _480_ (.I(_201_),
    .ZN(_237_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _481_ (.A1(\pll_control.tint[4] ),
    .A2(_190_),
    .A3(\pll_control.tint[1] ),
    .A4(_119_),
    .ZN(_238_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _482_ (.I(_191_),
    .ZN(_239_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _483_ (.A1(_121_),
    .A2(_202_),
    .B(_238_),
    .C(_239_),
    .ZN(_240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input27 (.I(ext_trim[3]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _485_ (.A1(net2),
    .A2(net14),
    .ZN(_242_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _486_ (.A1(_236_),
    .A2(_237_),
    .A3(_240_),
    .B(_242_),
    .ZN(\itrim[14] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _487_ (.A1(_230_),
    .A2(_200_),
    .A3(_212_),
    .ZN(_243_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _488_ (.I(_187_),
    .ZN(_244_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _489_ (.A1(_232_),
    .A2(_244_),
    .A3(_193_),
    .Z(_245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _490_ (.A1(net2),
    .A2(net15),
    .ZN(_246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _491_ (.A1(_243_),
    .A2(_245_),
    .B(_246_),
    .ZN(\itrim[15] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _492_ (.A1(_114_),
    .A2(_120_),
    .Z(_247_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _493_ (.A1(_247_),
    .A2(_115_),
    .A3(net2),
    .Z(_248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _494_ (.A1(net2),
    .A2(net16),
    .ZN(_249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _495_ (.A1(_248_),
    .A2(_249_),
    .ZN(\itrim[16] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _496_ (.A1(_236_),
    .A2(_213_),
    .ZN(_250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _497_ (.A1(_250_),
    .A2(_238_),
    .ZN(_251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _498_ (.A1(net2),
    .A2(net17),
    .ZN(_252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _499_ (.A1(_251_),
    .A2(_252_),
    .ZN(\itrim[17] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _500_ (.I(_194_),
    .ZN(_253_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _501_ (.A1(_188_),
    .A2(_231_),
    .A3(_253_),
    .Z(_254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _502_ (.A1(net2),
    .A2(net18),
    .ZN(_255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _503_ (.A1(_243_),
    .A2(_254_),
    .B(_255_),
    .ZN(\itrim[18] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _504_ (.A1(_226_),
    .A2(_115_),
    .ZN(_256_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _505_ (.I0(_256_),
    .I1(net19),
    .S(net2),
    .Z(\itrim[19] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _506_ (.A1(_239_),
    .A2(_202_),
    .B(\pll_control.tint[4] ),
    .ZN(_257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _507_ (.A1(net2),
    .A2(net20),
    .ZN(_258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _508_ (.A1(_237_),
    .A2(_257_),
    .B(_258_),
    .ZN(\itrim[1] ));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _509_ (.A1(\pll_control.tint[1] ),
    .A2(\pll_control.tint[2] ),
    .B(\pll_control.tint[3] ),
    .C(\pll_control.tint[4] ),
    .ZN(_259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _510_ (.A1(net2),
    .A2(net21),
    .ZN(_260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _511_ (.A1(_259_),
    .A2(net2),
    .B(_260_),
    .ZN(\itrim[20] ));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _512_ (.A1(_224_),
    .A2(_118_),
    .A3(\pll_control.tint[0] ),
    .Z(_261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _513_ (.A1(net2),
    .A2(net22),
    .ZN(_262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _514_ (.A1(_248_),
    .A2(_261_),
    .B(_262_),
    .ZN(\itrim[21] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _515_ (.A1(net2),
    .A2(net23),
    .Z(_263_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _516_ (.A1(_250_),
    .A2(_263_),
    .Z(\itrim[22] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _517_ (.I0(\pll_control.tint[4] ),
    .I1(net24),
    .S(net2),
    .Z(\itrim[23] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _518_ (.I0(_129_),
    .I1(net25),
    .S(net2),
    .Z(\itrim[24] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _519_ (.A1(net2),
    .A2(net26),
    .ZN(_264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _520_ (.A1(_243_),
    .A2(_195_),
    .B(_264_),
    .ZN(\itrim[25] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _521_ (.A1(_112_),
    .A2(_115_),
    .ZN(_265_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _522_ (.I0(_265_),
    .I1(net27),
    .S(net2),
    .Z(\itrim[2] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _523_ (.A1(net2),
    .A2(net28),
    .ZN(_266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _524_ (.A1(_244_),
    .A2(_266_),
    .ZN(\itrim[3] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _525_ (.A1(net2),
    .A2(net29),
    .ZN(_267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _526_ (.A1(_207_),
    .A2(_267_),
    .ZN(\itrim[4] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _527_ (.A1(net2),
    .A2(net30),
    .ZN(_268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _528_ (.A1(_237_),
    .A2(_268_),
    .ZN(\itrim[5] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _529_ (.A1(_182_),
    .A2(_118_),
    .ZN(_269_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _530_ (.I0(_269_),
    .I1(net31),
    .S(net2),
    .Z(\itrim[6] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _531_ (.A1(net2),
    .A2(net32),
    .ZN(_270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _532_ (.A1(_220_),
    .A2(_270_),
    .ZN(\itrim[7] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _533_ (.A1(net2),
    .A2(net33),
    .ZN(_271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _534_ (.A1(_195_),
    .A2(_271_),
    .ZN(\itrim[8] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _535_ (.A1(net2),
    .A2(net34),
    .ZN(_272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _536_ (.A1(_213_),
    .A2(_272_),
    .ZN(\itrim[9] ));
 gf180mcu_fd_sc_mcu7t5v0__addf_2 _537_ (.A(_000_),
    .B(\pll_control.count1[1] ),
    .CI(\pll_control.count0[1] ),
    .CO(_001_),
    .S(_273_));
 gf180mcu_fd_sc_mcu7t5v0__addf_2 _538_ (.A(_002_),
    .B(\pll_control.tval[0] ),
    .CI(\pll_control.tval[1] ),
    .CO(_003_),
    .S(_004_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _539_ (.A(\pll_control.count1[4] ),
    .B(\pll_control.count0[4] ),
    .CO(_005_),
    .S(_006_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _540_ (.A(\pll_control.count1[3] ),
    .B(\pll_control.count0[3] ),
    .CO(_007_),
    .S(_008_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _541_ (.A(\pll_control.count1[2] ),
    .B(\pll_control.count0[2] ),
    .CO(_009_),
    .S(_010_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _542_ (.A(\pll_control.count1[1] ),
    .B(\pll_control.count0[1] ),
    .CO(_011_),
    .S(_012_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _543_ (.A(_013_),
    .B(_014_),
    .CO(_015_),
    .S(_016_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _544_ (.A(_017_),
    .B(_018_),
    .CO(_019_),
    .S(_020_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _545_ (.A(_021_),
    .B(_022_),
    .CO(_023_),
    .S(_024_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _546_ (.A(_025_),
    .B(_273_),
    .CO(_026_),
    .S(_027_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _547_ (.A(\pll_control.count1[0] ),
    .B(\pll_control.count0[0] ),
    .CO(_000_),
    .S(_028_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _548_ (.A(net3),
    .B(_029_),
    .CO(_030_),
    .S(_031_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _549_ (.A(\pll_control.count0[0] ),
    .B(\pll_control.count0[1] ),
    .CO(_032_),
    .S(_033_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _550_ (.A(\pll_control.count0[4] ),
    .B(_034_),
    .CO(_035_),
    .S(_036_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _551_ (.A(_002_),
    .B(\pll_control.tval[1] ),
    .CO(_037_),
    .S(_038_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _552_ (.A(_002_),
    .B(\pll_control.tint[0] ),
    .CO(_039_),
    .S(_040_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _553_ (.A(_002_),
    .B(\pll_control.tint[1] ),
    .CO(_041_),
    .S(_042_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _554_ (.A(_002_),
    .B(\pll_control.tint[2] ),
    .CO(_043_),
    .S(_044_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _555_ (.A(_002_),
    .B(\pll_control.tint[3] ),
    .CO(_045_),
    .S(_046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input26 (.I(ext_trim[2]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count0[0]$_DFFE_PP0P_  (.D(_048_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.count0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count0[1]$_DFFE_PP0P_  (.D(_049_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.count0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count0[2]$_DFFE_PP0P_  (.D(_050_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.count0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count0[3]$_DFFE_PP0P_  (.D(_051_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.count0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count0[4]$_DFFE_PP0P_  (.D(_052_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.count0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count1[0]$_DFFE_PP0N_  (.D(_053_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.count1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count1[1]$_DFFE_PP0N_  (.D(_054_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.count1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count1[2]$_DFFE_PP0N_  (.D(_055_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.count1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count1[3]$_DFFE_PP0N_  (.D(_056_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.count1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.count1[4]$_DFFE_PP0N_  (.D(_057_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.count1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.oscbuf[0]$_DFF_PP0_  (.D(osc),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.oscbuf[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.oscbuf[1]$_DFF_PP0_  (.D(\pll_control.oscbuf[0] ),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.oscbuf[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.oscbuf[2]$_DFF_PP0_  (.D(\pll_control.oscbuf[1] ),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.oscbuf[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.prep[0]$_DFFE_PP0N_  (.D(_058_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.prep[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.prep[1]$_DFFE_PP0N_  (.D(_059_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.prep[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.prep[2]$_DFFE_PP0N_  (.D(_060_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.prep[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.tval[0]$_DFFE_PP0P_  (.D(_061_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.tval[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.tval[1]$_DFFE_PP0P_  (.D(_062_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.tval[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.tval[2]$_DFFE_PP0P_  (.D(_063_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.tint[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.tval[3]$_DFFE_PP0P_  (.D(_064_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.tint[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.tval[4]$_DFFE_PP0P_  (.D(_065_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.tint[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.tval[5]$_DFFE_PP0P_  (.D(_066_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.tint[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \pll_control.tval[6]$_DFFE_PP0P_  (.D(_067_),
    .RN(_047_),
    .CLK(net36),
    .Q(\pll_control.tint[4] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input25 (.I(ext_trim[25]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input24 (.I(ext_trim[24]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[0].id.delayen0  (.EN(\itrim[0] ),
    .I(\ringosc.dstage[0].id.d2 ),
    .ZN(\ringosc.dstage[0].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[0].id.delayen1  (.EN(\itrim[13] ),
    .I(\ringosc.dstage[0].id.in ),
    .ZN(\ringosc.dstage[0].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[0].id.delayenb0  (.EN(\ringosc.dstage[0].id.trim0b ),
    .I(\ringosc.dstage[0].id.in ),
    .ZN(\ringosc.dstage[0].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[0].id.delayenb1  (.EN(\ringosc.dstage[0].id.trim1b ),
    .I(\ringosc.dstage[0].id.in ),
    .ZN(\ringosc.dstage[0].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[0].id.delayint0  (.I(\ringosc.dstage[0].id.d1 ),
    .ZN(\ringosc.dstage[0].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[0].id.trim0bar  (.I(\itrim[0] ),
    .ZN(\ringosc.dstage[0].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[0].id.trim1bar  (.I(\itrim[13] ),
    .ZN(\ringosc.dstage[0].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input23 (.I(ext_trim[23]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input22 (.I(ext_trim[22]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[10].id.delayen0  (.EN(\itrim[10] ),
    .I(\ringosc.dstage[10].id.d2 ),
    .ZN(\ringosc.dstage[10].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[10].id.delayen1  (.EN(\itrim[23] ),
    .I(\ringosc.dstage[10].id.in ),
    .ZN(\ringosc.dstage[10].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[10].id.delayenb0  (.EN(\ringosc.dstage[10].id.trim0b ),
    .I(\ringosc.dstage[10].id.in ),
    .ZN(\ringosc.dstage[10].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[10].id.delayenb1  (.EN(\ringosc.dstage[10].id.trim1b ),
    .I(\ringosc.dstage[10].id.in ),
    .ZN(\ringosc.dstage[10].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[10].id.delayint0  (.I(\ringosc.dstage[10].id.d1 ),
    .ZN(\ringosc.dstage[10].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[10].id.trim0bar  (.I(\itrim[10] ),
    .ZN(\ringosc.dstage[10].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[10].id.trim1bar  (.I(\itrim[23] ),
    .ZN(\ringosc.dstage[10].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input21 (.I(ext_trim[21]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input20 (.I(ext_trim[20]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[11].id.delayen0  (.EN(\itrim[11] ),
    .I(\ringosc.dstage[11].id.d2 ),
    .ZN(\ringosc.dstage[11].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[11].id.delayen1  (.EN(\itrim[24] ),
    .I(\ringosc.dstage[10].id.out ),
    .ZN(\ringosc.dstage[11].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[11].id.delayenb0  (.EN(\ringosc.dstage[11].id.trim0b ),
    .I(\ringosc.dstage[10].id.out ),
    .ZN(\ringosc.dstage[11].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[11].id.delayenb1  (.EN(\ringosc.dstage[11].id.trim1b ),
    .I(\ringosc.dstage[10].id.out ),
    .ZN(\ringosc.dstage[11].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[11].id.delayint0  (.I(\ringosc.dstage[11].id.d1 ),
    .ZN(\ringosc.dstage[11].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[11].id.trim0bar  (.I(\itrim[11] ),
    .ZN(\ringosc.dstage[11].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[11].id.trim1bar  (.I(\itrim[24] ),
    .ZN(\ringosc.dstage[11].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input19 (.I(ext_trim[1]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input18 (.I(ext_trim[19]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[1].id.delayen0  (.EN(\itrim[1] ),
    .I(\ringosc.dstage[1].id.d2 ),
    .ZN(\ringosc.dstage[1].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[1].id.delayen1  (.EN(\itrim[14] ),
    .I(\ringosc.dstage[0].id.out ),
    .ZN(\ringosc.dstage[1].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[1].id.delayenb0  (.EN(\ringosc.dstage[1].id.trim0b ),
    .I(\ringosc.dstage[0].id.out ),
    .ZN(\ringosc.dstage[1].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[1].id.delayenb1  (.EN(\ringosc.dstage[1].id.trim1b ),
    .I(\ringosc.dstage[0].id.out ),
    .ZN(\ringosc.dstage[1].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[1].id.delayint0  (.I(\ringosc.dstage[1].id.d1 ),
    .ZN(\ringosc.dstage[1].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[1].id.trim0bar  (.I(\itrim[1] ),
    .ZN(\ringosc.dstage[1].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[1].id.trim1bar  (.I(\itrim[14] ),
    .ZN(\ringosc.dstage[1].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input17 (.I(ext_trim[18]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input16 (.I(ext_trim[17]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[2].id.delayen0  (.EN(\itrim[2] ),
    .I(\ringosc.dstage[2].id.d2 ),
    .ZN(\ringosc.dstage[2].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[2].id.delayen1  (.EN(\itrim[15] ),
    .I(\ringosc.dstage[1].id.out ),
    .ZN(\ringosc.dstage[2].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[2].id.delayenb0  (.EN(\ringosc.dstage[2].id.trim0b ),
    .I(\ringosc.dstage[1].id.out ),
    .ZN(\ringosc.dstage[2].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[2].id.delayenb1  (.EN(\ringosc.dstage[2].id.trim1b ),
    .I(\ringosc.dstage[1].id.out ),
    .ZN(\ringosc.dstage[2].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[2].id.delayint0  (.I(\ringosc.dstage[2].id.d1 ),
    .ZN(\ringosc.dstage[2].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[2].id.trim0bar  (.I(\itrim[2] ),
    .ZN(\ringosc.dstage[2].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[2].id.trim1bar  (.I(\itrim[15] ),
    .ZN(\ringosc.dstage[2].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input15 (.I(ext_trim[16]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input14 (.I(ext_trim[15]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[3].id.delayen0  (.EN(\itrim[3] ),
    .I(\ringosc.dstage[3].id.d2 ),
    .ZN(\ringosc.dstage[3].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[3].id.delayen1  (.EN(\itrim[16] ),
    .I(\ringosc.dstage[2].id.out ),
    .ZN(\ringosc.dstage[3].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[3].id.delayenb0  (.EN(\ringosc.dstage[3].id.trim0b ),
    .I(\ringosc.dstage[2].id.out ),
    .ZN(\ringosc.dstage[3].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[3].id.delayenb1  (.EN(\ringosc.dstage[3].id.trim1b ),
    .I(\ringosc.dstage[2].id.out ),
    .ZN(\ringosc.dstage[3].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[3].id.delayint0  (.I(\ringosc.dstage[3].id.d1 ),
    .ZN(\ringosc.dstage[3].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[3].id.trim0bar  (.I(\itrim[3] ),
    .ZN(\ringosc.dstage[3].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[3].id.trim1bar  (.I(\itrim[16] ),
    .ZN(\ringosc.dstage[3].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input13 (.I(ext_trim[14]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input12 (.I(ext_trim[13]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[4].id.delayen0  (.EN(\itrim[4] ),
    .I(\ringosc.dstage[4].id.d2 ),
    .ZN(\ringosc.dstage[4].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[4].id.delayen1  (.EN(\itrim[17] ),
    .I(\ringosc.dstage[3].id.out ),
    .ZN(\ringosc.dstage[4].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[4].id.delayenb0  (.EN(\ringosc.dstage[4].id.trim0b ),
    .I(\ringosc.dstage[3].id.out ),
    .ZN(\ringosc.dstage[4].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[4].id.delayenb1  (.EN(\ringosc.dstage[4].id.trim1b ),
    .I(\ringosc.dstage[3].id.out ),
    .ZN(\ringosc.dstage[4].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[4].id.delayint0  (.I(\ringosc.dstage[4].id.d1 ),
    .ZN(\ringosc.dstage[4].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[4].id.trim0bar  (.I(\itrim[4] ),
    .ZN(\ringosc.dstage[4].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[4].id.trim1bar  (.I(\itrim[17] ),
    .ZN(\ringosc.dstage[4].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input11 (.I(ext_trim[12]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input10 (.I(ext_trim[11]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[5].id.delayen0  (.EN(\itrim[5] ),
    .I(\ringosc.dstage[5].id.d2 ),
    .ZN(\ringosc.dstage[5].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[5].id.delayen1  (.EN(\itrim[18] ),
    .I(\ringosc.dstage[4].id.out ),
    .ZN(\ringosc.dstage[5].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[5].id.delayenb0  (.EN(\ringosc.dstage[5].id.trim0b ),
    .I(\ringosc.dstage[4].id.out ),
    .ZN(\ringosc.dstage[5].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[5].id.delayenb1  (.EN(\ringosc.dstage[5].id.trim1b ),
    .I(\ringosc.dstage[4].id.out ),
    .ZN(\ringosc.dstage[5].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[5].id.delayint0  (.I(\ringosc.dstage[5].id.d1 ),
    .ZN(\ringosc.dstage[5].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[5].id.trim0bar  (.I(\itrim[5] ),
    .ZN(\ringosc.dstage[5].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[5].id.trim1bar  (.I(\itrim[18] ),
    .ZN(\ringosc.dstage[5].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input9 (.I(ext_trim[10]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input8 (.I(ext_trim[0]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[6].id.delayen0  (.EN(\itrim[6] ),
    .I(\ringosc.dstage[6].id.d2 ),
    .ZN(\ringosc.dstage[6].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[6].id.delayen1  (.EN(\itrim[19] ),
    .I(\ringosc.dstage[5].id.out ),
    .ZN(\ringosc.dstage[6].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[6].id.delayenb0  (.EN(\ringosc.dstage[6].id.trim0b ),
    .I(\ringosc.dstage[5].id.out ),
    .ZN(\ringosc.dstage[6].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[6].id.delayenb1  (.EN(\ringosc.dstage[6].id.trim1b ),
    .I(\ringosc.dstage[5].id.out ),
    .ZN(\ringosc.dstage[6].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[6].id.delayint0  (.I(\ringosc.dstage[6].id.d1 ),
    .ZN(\ringosc.dstage[6].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[6].id.trim0bar  (.I(\itrim[6] ),
    .ZN(\ringosc.dstage[6].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[6].id.trim1bar  (.I(\itrim[19] ),
    .ZN(\ringosc.dstage[6].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input7 (.I(enable),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input6 (.I(div[4]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[7].id.delayen0  (.EN(\itrim[7] ),
    .I(\ringosc.dstage[7].id.d2 ),
    .ZN(\ringosc.dstage[7].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[7].id.delayen1  (.EN(\itrim[20] ),
    .I(\ringosc.dstage[6].id.out ),
    .ZN(\ringosc.dstage[7].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[7].id.delayenb0  (.EN(\ringosc.dstage[7].id.trim0b ),
    .I(\ringosc.dstage[6].id.out ),
    .ZN(\ringosc.dstage[7].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[7].id.delayenb1  (.EN(\ringosc.dstage[7].id.trim1b ),
    .I(\ringosc.dstage[6].id.out ),
    .ZN(\ringosc.dstage[7].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[7].id.delayint0  (.I(\ringosc.dstage[7].id.d1 ),
    .ZN(\ringosc.dstage[7].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[7].id.trim0bar  (.I(\itrim[7] ),
    .ZN(\ringosc.dstage[7].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[7].id.trim1bar  (.I(\itrim[20] ),
    .ZN(\ringosc.dstage[7].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input5 (.I(div[3]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input4 (.I(div[2]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[8].id.delayen0  (.EN(\itrim[8] ),
    .I(\ringosc.dstage[8].id.d2 ),
    .ZN(\ringosc.dstage[8].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[8].id.delayen1  (.EN(\itrim[21] ),
    .I(\ringosc.dstage[7].id.out ),
    .ZN(\ringosc.dstage[8].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[8].id.delayenb0  (.EN(\ringosc.dstage[8].id.trim0b ),
    .I(\ringosc.dstage[7].id.out ),
    .ZN(\ringosc.dstage[8].id.out ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[8].id.delayenb1  (.EN(\ringosc.dstage[8].id.trim1b ),
    .I(\ringosc.dstage[7].id.out ),
    .ZN(\ringosc.dstage[8].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[8].id.delayint0  (.I(\ringosc.dstage[8].id.d1 ),
    .ZN(\ringosc.dstage[8].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[8].id.trim0bar  (.I(\itrim[8] ),
    .ZN(\ringosc.dstage[8].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[8].id.trim1bar  (.I(\itrim[21] ),
    .ZN(\ringosc.dstage[8].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input3 (.I(div[1]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input2 (.I(div[0]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[9].id.delayen0  (.EN(\itrim[9] ),
    .I(\ringosc.dstage[9].id.d2 ),
    .ZN(\ringosc.dstage[10].id.in ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[9].id.delayen1  (.EN(\itrim[22] ),
    .I(\ringosc.dstage[8].id.out ),
    .ZN(\ringosc.dstage[9].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.dstage[9].id.delayenb0  (.EN(\ringosc.dstage[9].id.trim0b ),
    .I(\ringosc.dstage[8].id.out ),
    .ZN(\ringosc.dstage[10].id.in ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.dstage[9].id.delayenb1  (.EN(\ringosc.dstage[9].id.trim1b ),
    .I(\ringosc.dstage[8].id.out ),
    .ZN(\ringosc.dstage[9].id.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[9].id.delayint0  (.I(\ringosc.dstage[9].id.d1 ),
    .ZN(\ringosc.dstage[9].id.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[9].id.trim0bar  (.I(\itrim[9] ),
    .ZN(\ringosc.dstage[9].id.trim0b ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.dstage[9].id.trim1bar  (.I(\itrim[22] ),
    .ZN(\ringosc.dstage[9].id.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 \ringosc.ibufp00  (.I(\ringosc.dstage[0].id.in ),
    .ZN(\ringosc.c[0] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_12 \ringosc.ibufp01  (.I(\ringosc.c[0] ),
    .ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.ibufp10  (.I(\ringosc.dstage[5].id.out ),
    .ZN(\ringosc.c[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.ibufp11  (.I(\ringosc.c[1] ),
    .ZN(net37));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 \ringosc.iss.ctrlen0  (.A1(ireset),
    .A2(\itrim[12] ),
    .ZN(\ringosc.iss.ctrl0b ));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 input1 (.I(dco),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.iss.delayen0  (.EN(\itrim[12] ),
    .I(\ringosc.iss.d2 ),
    .ZN(\ringosc.dstage[0].id.in ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.iss.delayen1  (.EN(\itrim[25] ),
    .I(\ringosc.dstage[11].id.out ),
    .ZN(\ringosc.iss.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.iss.delayenb0  (.EN(\ringosc.iss.ctrl0b ),
    .I(\ringosc.dstage[11].id.out ),
    .ZN(\ringosc.dstage[0].id.in ));
 gf180mcu_fd_sc_mcu7t5v0__invz_2 \ringosc.iss.delayenb1  (.EN(\ringosc.iss.trim1b ),
    .I(\ringosc.dstage[11].id.out ),
    .ZN(\ringosc.iss.d1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.iss.delayint0  (.I(\ringosc.iss.d1 ),
    .ZN(\ringosc.iss.d2 ));
 gf180mcu_fd_sc_mcu7t5v0__invz_16 \ringosc.iss.reseten0  (.EN(ireset),
    .I(net1),
    .ZN(\ringosc.dstage[0].id.in ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \ringosc.iss.trim1bar  (.I(\itrim[25] ),
    .ZN(\ringosc.iss.trim1b ));
 gf180mcu_fd_sc_mcu7t5v0__tieh \ringosc.iss.reseten0_1  (.Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_193 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input33 (.I(ext_trim[9]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input34 (.I(resetb),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output35 (.I(net36),
    .Z(clockp[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output36 (.I(net37),
    .Z(clockp[1]));
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_0_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_0_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_0_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_0_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_0_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_0_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_0_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_0_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_1_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_1_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_1_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_1_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_1_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_1_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_1_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_2_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_2_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_2_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_2_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_2_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_2_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_2_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_2_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_2_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_3_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_3_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_3_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_3_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_3_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_3_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_4_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_4_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_4_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_4_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_4_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_4_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_5_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_5_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_5_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_5_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_5_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_5_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_5_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_5_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_5_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_6_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_6_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_6_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_6_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_6_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_6_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_7_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_7_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_7_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_7_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_8_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_8_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_8_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_8_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_8_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_8_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_9_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_9_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_9_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_9_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_9_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_9_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_9_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_10_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_10_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_10_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_10_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_10_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_10_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_10_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_10_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_10_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_11_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_11_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_11_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_11_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_11_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_11_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_11_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_11_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_11_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_11_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_11_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_12_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_12_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_12_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_12_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_12_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_12_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_12_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_12_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_12_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_12_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_12_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_13_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_13_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_13_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_13_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_13_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_13_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_13_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_13_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_13_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_13_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_14_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_14_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_14_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_14_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_14_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_14_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_14_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_14_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_14_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_15_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_15_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_15_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_15_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_15_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_15_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_15_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_15_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_15_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_15_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_16_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_16_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_16_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_16_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_16_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_16_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_16_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_16_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_16_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_16_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_16_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_16_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_16_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_16_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_17_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_17_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_17_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_17_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_17_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_17_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_17_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_17_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_18_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_18_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_18_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_18_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_18_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_18_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_19_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_19_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_19_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_19_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_19_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_19_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_19_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_19_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_19_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_20_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_20_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_20_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_20_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_20_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_20_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_20_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_20_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_20_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_20_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_20_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_20_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_21_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_21_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_21_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_21_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_21_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_21_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_21_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_21_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_22_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_22_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_22_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_22_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_22_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_22_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_22_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_22_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_22_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_23_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_23_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_23_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_23_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_23_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_23_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_23_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_23_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_23_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_23_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_23_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_23_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_23_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_23_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_23_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_23_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_23_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_23_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_24_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_24_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_24_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_24_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_24_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_24_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_24_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_24_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_25_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_25_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_25_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_25_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_25_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_25_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_25_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_25_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_25_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_26_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_26_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_26_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_26_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_26_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_26_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_26_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_26_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_26_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_26_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_26_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_27_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_27_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_27_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_27_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_27_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_27_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_27_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_27_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_27_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_27_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_27_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_27_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_28_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_28_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_28_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_28_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_28_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_28_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_28_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_28_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_28_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_28_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_28_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_29_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_29_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_29_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_29_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_29_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_29_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_29_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_29_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_29_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_29_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_29_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_29_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_29_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_29_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_30_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_30_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_30_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_30_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_30_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_30_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_30_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_30_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_30_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_30_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_31_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_31_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_31_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_31_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_31_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_31_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_31_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_31_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_31_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_31_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_31_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_31_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_31_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_32_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_32_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_32_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_32_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_32_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_32_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_32_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_32_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_32_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_32_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_33_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_33_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_33_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_33_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_33_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_33_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_33_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_33_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_33_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_33_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_33_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_33_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_34_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_34_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_34_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_34_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_34_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_34_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_34_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_34_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_34_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_34_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_34_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_35_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_35_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_35_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_35_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_35_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_35_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_35_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_35_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_35_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_35_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_35_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_36_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_36_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_36_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_36_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_36_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_36_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_36_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_36_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_36_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_36_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_36_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_36_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_36_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_36_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_36_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_37_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_37_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_37_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_37_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_37_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_37_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_37_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_37_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_37_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_37_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_37_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_37_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_37_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_38_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_38_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_38_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_38_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_38_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_38_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_38_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_38_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_38_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_38_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_38_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_39_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_39_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_39_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_39_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_39_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_39_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_39_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_39_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_39_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_40_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_40_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_40_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_40_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_40_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_40_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_40_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_40_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_40_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_40_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_41_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_41_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_41_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_41_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_41_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_41_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_41_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_41_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_41_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_41_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_42_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_42_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_42_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_42_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_42_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_42_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_42_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_42_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_42_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_42_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_42_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_42_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_42_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_43_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_43_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_43_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_43_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_43_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_43_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_43_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_43_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_43_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_43_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_43_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_44_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_44_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_44_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_44_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_44_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_44_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_44_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_44_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_44_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_45_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_45_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_45_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_45_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_45_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_45_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_45_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_45_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_45_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_45_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_45_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_45_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_46_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_46_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_46_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_46_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_46_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_46_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_46_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_46_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_46_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_46_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_46_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_47_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_47_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_47_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_47_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_47_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_47_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_47_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_48_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_48_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_48_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_48_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_48_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_48_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_49_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_49_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_49_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_49_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_49_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_49_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_49_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_49_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_49_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_49_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_50_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_50_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_50_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_50_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_50_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_50_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_50_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_50_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_51_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_51_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_51_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_51_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_51_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_51_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_51_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_52_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_52_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_52_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_52_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_52_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_52_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_52_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_53_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_53_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_53_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_53_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_53_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_53_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_53_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_53_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_53_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_53_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_53_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_53_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_53_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_53_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_54_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_54_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_54_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_54_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_54_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_54_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_54_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_55_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_55_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_55_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_55_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_55_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_55_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_55_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_56_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_56_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_56_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_56_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_56_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_56_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_56_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_56_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_56_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_56_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_56_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_57_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_57_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_57_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_57_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_57_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_57_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_57_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_57_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_57_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_57_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_57_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_57_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_58_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_58_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_58_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_58_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_58_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_58_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_58_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_58_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_59_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_59_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_59_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_59_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_59_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_59_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_60_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_60_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_60_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_60_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_60_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_60_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_60_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_60_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_60_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_60_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_60_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_60_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_61_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_61_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_61_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_61_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_61_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_61_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_61_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_61_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_61_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_61_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_62_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_62_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_62_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_62_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_62_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_62_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_62_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_62_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_63_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_63_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_63_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_63_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_63_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_63_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_63_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_448 ();
endmodule
