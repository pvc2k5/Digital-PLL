VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

VIA ring_osc2x13_via1_2_8960_1800_1_4_1240_1240
  VIARULE Via1_GEN_HH ;
  CUTSIZE 0.26 0.26 ;
  LAYERS Metal1 Via1 Metal2 ;
  CUTSPACING 0.36 0.36 ;
  ENCLOSURE 0.06 0.32 0.01 0.06 ;
  ROWCOL 1 4 ;
END ring_osc2x13_via1_2_8960_1800_1_4_1240_1240

VIA ring_osc2x13_via2_3_8960_560_1_8_1040_1040
  VIARULE Via2_GEN_HH ;
  CUTSIZE 0.26 0.26 ;
  LAYERS Metal2 Via2 Metal3 ;
  CUTSPACING 0.26 0.26 ;
  ENCLOSURE 0.01 0.06 0.06 0.01 ;
  ROWCOL 1 8 ;
END ring_osc2x13_via2_3_8960_560_1_8_1040_1040

VIA ring_osc2x13_via3_4_8960_560_1_8_1040_1040
  VIARULE Via3_GEN_HH ;
  CUTSIZE 0.26 0.26 ;
  LAYERS Metal3 Via3 Metal4 ;
  CUTSPACING 0.26 0.26 ;
  ENCLOSURE 0.06 0.01 0.29 0.06 ;
  ROWCOL 1 8 ;
END ring_osc2x13_via3_4_8960_560_1_8_1040_1040

MACRO ring_osc2x13
  FOREIGN ring_osc2x13 0 0 ;
  CLASS BLOCK ;
  SIZE 142.64 BY 142.64 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER Metal4 ;
        RECT  117.04 7.39 121.52 133.73 ;
        RECT  72.24 7.39 76.72 133.73 ;
        RECT  27.44 7.39 31.92 133.73 ;
      LAYER Metal1 ;
        RECT  2.24 132.83 140.56 133.73 ;
        RECT  2.24 124.99 140.56 125.89 ;
        RECT  2.24 117.15 140.56 118.05 ;
        RECT  2.24 109.31 140.56 110.21 ;
        RECT  2.24 101.47 140.56 102.37 ;
        RECT  2.24 93.63 140.56 94.53 ;
        RECT  2.24 85.79 140.56 86.69 ;
        RECT  2.24 77.95 140.56 78.85 ;
        RECT  2.24 70.11 140.56 71.01 ;
        RECT  2.24 62.27 140.56 63.17 ;
        RECT  2.24 54.43 140.56 55.33 ;
        RECT  2.24 46.59 140.56 47.49 ;
        RECT  2.24 38.75 140.56 39.65 ;
        RECT  2.24 30.91 140.56 31.81 ;
        RECT  2.24 23.07 140.56 23.97 ;
        RECT  2.24 15.23 140.56 16.13 ;
        RECT  2.24 7.39 140.56 8.29 ;
      VIA 119.28 133.28 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 133.28 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 133.28 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 125.44 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 125.44 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 125.44 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 117.6 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 117.6 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 117.6 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 109.76 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 109.76 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 109.76 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 101.92 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 101.92 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 101.92 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 94.08 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 94.08 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 94.08 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 86.24 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 86.24 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 86.24 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 78.4 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 78.4 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 78.4 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 70.56 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 70.56 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 70.56 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 62.72 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 62.72 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 62.72 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 54.88 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 54.88 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 54.88 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 47.04 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 47.04 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 47.04 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 39.2 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 39.2 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 39.2 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 31.36 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 31.36 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 31.36 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 23.52 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 23.52 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 23.52 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 15.68 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 15.68 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 15.68 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 119.28 7.84 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 119.28 7.84 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 119.28 7.84 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 133.28 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 133.28 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 133.28 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 125.44 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 125.44 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 125.44 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 117.6 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 117.6 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 117.6 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 109.76 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 109.76 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 109.76 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 101.92 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 101.92 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 101.92 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 94.08 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 94.08 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 94.08 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 86.24 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 86.24 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 86.24 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 78.4 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 78.4 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 78.4 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 70.56 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 70.56 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 70.56 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 62.72 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 62.72 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 62.72 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 54.88 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 54.88 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 54.88 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 47.04 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 47.04 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 47.04 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 39.2 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 39.2 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 39.2 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 31.36 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 31.36 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 31.36 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 23.52 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 23.52 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 23.52 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 15.68 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 15.68 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 15.68 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 74.48 7.84 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 74.48 7.84 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 74.48 7.84 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 133.28 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 133.28 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 133.28 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 125.44 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 125.44 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 125.44 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 117.6 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 117.6 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 117.6 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 109.76 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 109.76 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 109.76 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 101.92 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 101.92 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 101.92 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 94.08 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 94.08 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 94.08 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 86.24 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 86.24 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 86.24 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 78.4 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 78.4 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 78.4 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 70.56 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 70.56 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 70.56 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 62.72 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 62.72 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 62.72 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 54.88 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 54.88 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 54.88 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 47.04 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 47.04 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 47.04 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 39.2 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 39.2 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 39.2 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 31.36 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 31.36 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 31.36 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 23.52 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 23.52 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 23.52 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 15.68 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 15.68 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 15.68 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 29.68 7.84 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 29.68 7.84 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 29.68 7.84 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER Metal4 ;
        RECT  112 3.47 116.48 137.65 ;
        RECT  67.2 3.47 71.68 137.65 ;
        RECT  22.4 3.47 26.88 137.65 ;
      LAYER Metal1 ;
        RECT  2.24 136.75 140.56 137.65 ;
        RECT  2.24 128.91 140.56 129.81 ;
        RECT  2.24 121.07 140.56 121.97 ;
        RECT  2.24 113.23 140.56 114.13 ;
        RECT  2.24 105.39 140.56 106.29 ;
        RECT  2.24 97.55 140.56 98.45 ;
        RECT  2.24 89.71 140.56 90.61 ;
        RECT  2.24 81.87 140.56 82.77 ;
        RECT  2.24 74.03 140.56 74.93 ;
        RECT  2.24 66.19 140.56 67.09 ;
        RECT  2.24 58.35 140.56 59.25 ;
        RECT  2.24 50.51 140.56 51.41 ;
        RECT  2.24 42.67 140.56 43.57 ;
        RECT  2.24 34.83 140.56 35.73 ;
        RECT  2.24 26.99 140.56 27.89 ;
        RECT  2.24 19.15 140.56 20.05 ;
        RECT  2.24 11.31 140.56 12.21 ;
        RECT  2.24 3.47 140.56 4.37 ;
      VIA 114.24 137.2 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 137.2 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 137.2 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 129.36 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 129.36 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 129.36 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 121.52 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 121.52 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 121.52 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 113.68 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 113.68 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 113.68 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 105.84 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 105.84 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 105.84 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 98 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 98 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 98 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 90.16 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 90.16 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 90.16 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 82.32 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 82.32 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 82.32 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 74.48 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 74.48 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 74.48 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 66.64 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 66.64 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 66.64 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 58.8 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 58.8 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 58.8 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 50.96 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 50.96 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 50.96 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 43.12 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 43.12 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 43.12 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 35.28 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 35.28 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 35.28 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 27.44 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 27.44 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 27.44 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 19.6 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 19.6 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 19.6 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 11.76 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 11.76 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 11.76 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 114.24 3.92 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 114.24 3.92 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 114.24 3.92 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 137.2 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 137.2 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 137.2 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 129.36 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 129.36 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 129.36 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 121.52 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 121.52 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 121.52 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 113.68 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 113.68 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 113.68 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 105.84 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 105.84 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 105.84 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 98 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 98 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 98 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 90.16 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 90.16 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 90.16 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 82.32 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 82.32 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 82.32 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 74.48 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 74.48 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 74.48 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 66.64 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 66.64 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 66.64 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 58.8 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 58.8 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 58.8 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 50.96 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 50.96 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 50.96 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 43.12 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 43.12 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 43.12 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 35.28 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 35.28 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 35.28 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 27.44 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 27.44 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 27.44 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 19.6 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 19.6 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 19.6 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 11.76 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 11.76 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 11.76 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 69.44 3.92 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 69.44 3.92 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 69.44 3.92 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 137.2 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 137.2 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 137.2 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 129.36 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 129.36 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 129.36 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 121.52 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 121.52 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 121.52 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 113.68 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 113.68 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 113.68 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 105.84 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 105.84 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 105.84 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 98 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 98 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 98 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 90.16 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 90.16 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 90.16 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 82.32 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 82.32 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 82.32 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 74.48 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 74.48 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 74.48 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 66.64 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 66.64 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 66.64 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 58.8 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 58.8 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 58.8 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 50.96 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 50.96 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 50.96 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 43.12 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 43.12 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 43.12 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 35.28 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 35.28 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 35.28 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 27.44 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 27.44 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 27.44 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 19.6 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 19.6 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 19.6 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 11.76 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 11.76 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 11.76 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
      VIA 24.64 3.92 ring_osc2x13_via3_4_8960_560_1_8_1040_1040 ;
      VIA 24.64 3.92 ring_osc2x13_via2_3_8960_560_1_8_1040_1040 ;
      VIA 24.64 3.92 ring_osc2x13_via1_2_8960_1800_1_4_1240_1240 ;
    END
  END VSS
  PIN clockp[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  128.1 142.12 128.38 142.64 ;
    END
  END clockp[0]
  PIN clockp[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  44.1 142.12 44.38 142.64 ;
    END
  END clockp[1]
  PIN dco
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  57.54 142.12 57.82 142.64 ;
    END
  END dco
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  100.1 142.12 100.38 142.64 ;
    END
  END enable
  PIN ext_trim[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  114.66 142.12 114.94 142.64 ;
    END
  END ext_trim[0]
  PIN ext_trim[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  78.82 142.12 79.1 142.64 ;
    END
  END ext_trim[10]
  PIN ext_trim[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  94.5 142.12 94.78 142.64 ;
    END
  END ext_trim[11]
  PIN ext_trim[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  101.22 142.12 101.5 142.64 ;
    END
  END ext_trim[12]
  PIN ext_trim[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  106.82 142.12 107.1 142.64 ;
    END
  END ext_trim[13]
  PIN ext_trim[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  90.02 142.12 90.3 142.64 ;
    END
  END ext_trim[14]
  PIN ext_trim[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  105.7 142.12 105.98 142.64 ;
    END
  END ext_trim[15]
  PIN ext_trim[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  79.94 142.12 80.22 142.64 ;
    END
  END ext_trim[16]
  PIN ext_trim[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  70.98 142.12 71.26 142.64 ;
    END
  END ext_trim[17]
  PIN ext_trim[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  66.5 142.12 66.78 142.64 ;
    END
  END ext_trim[18]
  PIN ext_trim[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  23.94 142.12 24.22 142.64 ;
    END
  END ext_trim[19]
  PIN ext_trim[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  87.78 142.12 88.06 142.64 ;
    END
  END ext_trim[1]
  PIN ext_trim[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  27.3 142.12 27.58 142.64 ;
    END
  END ext_trim[20]
  PIN ext_trim[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  28.42 142.12 28.7 142.64 ;
    END
  END ext_trim[21]
  PIN ext_trim[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  53.06 142.12 53.34 142.64 ;
    END
  END ext_trim[22]
  PIN ext_trim[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  72.1 142.12 72.38 142.64 ;
    END
  END ext_trim[23]
  PIN ext_trim[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  77.7 142.12 77.98 142.64 ;
    END
  END ext_trim[24]
  PIN ext_trim[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  113.54 142.12 113.82 142.64 ;
    END
  END ext_trim[25]
  PIN ext_trim[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  103.46 142.12 103.74 142.64 ;
    END
  END ext_trim[2]
  PIN ext_trim[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  73.22 142.12 73.5 142.64 ;
    END
  END ext_trim[3]
  PIN ext_trim[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  45.22 142.12 45.5 142.64 ;
    END
  END ext_trim[4]
  PIN ext_trim[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  47.46 142.12 47.74 142.64 ;
    END
  END ext_trim[5]
  PIN ext_trim[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  22.82 142.12 23.1 142.64 ;
    END
  END ext_trim[6]
  PIN ext_trim[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  21.7 142.12 21.98 142.64 ;
    END
  END ext_trim[7]
  PIN ext_trim[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  42.98 142.12 43.26 142.64 ;
    END
  END ext_trim[8]
  PIN ext_trim[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  55.3 142.12 55.58 142.64 ;
    END
  END ext_trim[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  102.34 142.12 102.62 142.64 ;
    END
  END reset
  PIN trim[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  112.42 142.12 112.7 142.64 ;
    END
  END trim[0]
  PIN trim[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  82.18 142.12 82.46 142.64 ;
    END
  END trim[10]
  PIN trim[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  97.86 142.12 98.14 142.64 ;
    END
  END trim[11]
  PIN trim[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  104.58 142.12 104.86 142.64 ;
    END
  END trim[12]
  PIN trim[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  110.18 142.12 110.46 142.64 ;
    END
  END trim[13]
  PIN trim[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  93.38 142.12 93.66 142.64 ;
    END
  END trim[14]
  PIN trim[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  109.06 142.12 109.34 142.64 ;
    END
  END trim[15]
  PIN trim[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  84.42 142.12 84.7 142.64 ;
    END
  END trim[16]
  PIN trim[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  74.34 142.12 74.62 142.64 ;
    END
  END trim[17]
  PIN trim[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  69.86 142.12 70.14 142.64 ;
    END
  END trim[18]
  PIN trim[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  29.54 142.12 29.82 142.64 ;
    END
  END trim[19]
  PIN trim[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  91.14 142.12 91.42 142.64 ;
    END
  END trim[1]
  PIN trim[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  30.66 142.12 30.94 142.64 ;
    END
  END trim[20]
  PIN trim[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  31.78 142.12 32.06 142.64 ;
    END
  END trim[21]
  PIN trim[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  56.42 142.12 56.7 142.64 ;
    END
  END trim[22]
  PIN trim[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  75.46 142.12 75.74 142.64 ;
    END
  END trim[23]
  PIN trim[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  81.06 142.12 81.34 142.64 ;
    END
  END trim[24]
  PIN trim[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  111.3 142.12 111.58 142.64 ;
    END
  END trim[25]
  PIN trim[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  107.94 142.12 108.22 142.64 ;
    END
  END trim[2]
  PIN trim[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  76.58 142.12 76.86 142.64 ;
    END
  END trim[3]
  PIN trim[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  48.58 142.12 48.86 142.64 ;
    END
  END trim[4]
  PIN trim[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  50.82 142.12 51.1 142.64 ;
    END
  END trim[5]
  PIN trim[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  26.18 142.12 26.46 142.64 ;
    END
  END trim[6]
  PIN trim[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  25.06 142.12 25.34 142.64 ;
    END
  END trim[7]
  PIN trim[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  46.34 142.12 46.62 142.64 ;
    END
  END trim[8]
  PIN trim[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT  58.66 142.12 58.94 142.64 ;
    END
  END trim[9]
  OBS
    LAYER Metal1 ;
     RECT  2.24 3.47 140.56 142.64 ;
    LAYER Metal2 ;
     RECT  2.24 3.47 140.56 142.64 ;
    LAYER Metal3 ;
     RECT  2.24 3.47 140.56 142.64 ;
    LAYER Metal4 ;
     RECT  2.24 3.47 140.56 142.64 ;
  END
END ring_osc2x13
END LIBRARY
